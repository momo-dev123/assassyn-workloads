VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA run_benchmark_via1_2_72630_18_1_2017_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 2017 ;
END run_benchmark_via1_2_72630_18_1_2017_36_36

VIA run_benchmark_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END run_benchmark_VIA23_1_3_36_36

VIA run_benchmark_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END run_benchmark_VIA34_1_2_58_52

VIA run_benchmark_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END run_benchmark_VIA45_1_2_58_58

VIA run_benchmark_via5_6_120_288_1_2_58_322
  VIARULE M6_M5widePWR1p152 ;
  CUTSIZE 0.024 0.288 ;
  LAYERS M5 V5 M6 ;
  CUTSPACING 0.034 0.034 ;
  ENCLOSURE 0.019 0 0 0 ;
  ROWCOL 1 2 ;
END run_benchmark_via5_6_120_288_1_2_58_322

MACRO run_benchmark
  FOREIGN run_benchmark 0 0 ;
  CLASS BLOCK ;
  SIZE 74.707 BY 74.707 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.458 67.833 72.426 68.121 ;
        RECT  1.458 61.833 72.426 62.121 ;
        RECT  1.458 55.833 72.426 56.121 ;
        RECT  1.458 49.833 72.426 50.121 ;
        RECT  1.458 43.833 72.426 44.121 ;
        RECT  1.458 37.833 72.426 38.121 ;
        RECT  1.458 31.833 72.426 32.121 ;
        RECT  1.458 25.833 72.426 26.121 ;
        RECT  1.458 19.833 72.426 20.121 ;
        RECT  1.458 13.833 72.426 14.121 ;
        RECT  1.458 7.833 72.426 8.121 ;
        RECT  1.458 1.833 72.426 2.121 ;
      LAYER M5 ;
        RECT  72.306 1.327 72.426 73.193 ;
        RECT  66.402 1.327 66.522 73.193 ;
        RECT  60.498 1.327 60.618 73.193 ;
        RECT  54.594 1.327 54.714 73.193 ;
        RECT  48.69 1.327 48.81 73.193 ;
        RECT  42.786 1.327 42.906 73.193 ;
        RECT  36.882 1.327 37.002 73.193 ;
        RECT  30.978 1.327 31.098 73.193 ;
        RECT  25.074 1.327 25.194 73.193 ;
        RECT  19.17 1.327 19.29 73.193 ;
        RECT  13.266 1.327 13.386 73.193 ;
        RECT  7.362 1.327 7.482 73.193 ;
        RECT  1.458 1.327 1.578 73.193 ;
      LAYER M2 ;
        RECT  1.026 73.161 73.656 73.179 ;
        RECT  1.026 72.621 73.656 72.639 ;
        RECT  1.026 72.081 73.656 72.099 ;
        RECT  1.026 71.541 73.656 71.559 ;
        RECT  1.026 71.001 73.656 71.019 ;
        RECT  1.026 70.461 73.656 70.479 ;
        RECT  1.026 69.921 73.656 69.939 ;
        RECT  1.026 69.381 73.656 69.399 ;
        RECT  1.026 68.841 73.656 68.859 ;
        RECT  1.026 68.301 73.656 68.319 ;
        RECT  1.026 67.761 73.656 67.779 ;
        RECT  1.026 67.221 73.656 67.239 ;
        RECT  1.026 66.681 73.656 66.699 ;
        RECT  1.026 66.141 73.656 66.159 ;
        RECT  1.026 65.601 73.656 65.619 ;
        RECT  1.026 65.061 73.656 65.079 ;
        RECT  1.026 64.521 73.656 64.539 ;
        RECT  1.026 63.981 73.656 63.999 ;
        RECT  1.026 63.441 73.656 63.459 ;
        RECT  1.026 62.901 73.656 62.919 ;
        RECT  1.026 62.361 73.656 62.379 ;
        RECT  1.026 61.821 73.656 61.839 ;
        RECT  1.026 61.281 73.656 61.299 ;
        RECT  1.026 60.741 73.656 60.759 ;
        RECT  1.026 60.201 73.656 60.219 ;
        RECT  1.026 59.661 73.656 59.679 ;
        RECT  1.026 59.121 73.656 59.139 ;
        RECT  1.026 58.581 73.656 58.599 ;
        RECT  1.026 58.041 73.656 58.059 ;
        RECT  1.026 57.501 73.656 57.519 ;
        RECT  1.026 56.961 73.656 56.979 ;
        RECT  1.026 56.421 73.656 56.439 ;
        RECT  1.026 55.881 73.656 55.899 ;
        RECT  1.026 55.341 73.656 55.359 ;
        RECT  1.026 54.801 73.656 54.819 ;
        RECT  1.026 54.261 73.656 54.279 ;
        RECT  1.026 53.721 73.656 53.739 ;
        RECT  1.026 53.181 73.656 53.199 ;
        RECT  1.026 52.641 73.656 52.659 ;
        RECT  1.026 52.101 73.656 52.119 ;
        RECT  1.026 51.561 73.656 51.579 ;
        RECT  1.026 51.021 73.656 51.039 ;
        RECT  1.026 50.481 73.656 50.499 ;
        RECT  1.026 49.941 73.656 49.959 ;
        RECT  1.026 49.401 73.656 49.419 ;
        RECT  1.026 48.861 73.656 48.879 ;
        RECT  1.026 48.321 73.656 48.339 ;
        RECT  1.026 47.781 73.656 47.799 ;
        RECT  1.026 47.241 73.656 47.259 ;
        RECT  1.026 46.701 73.656 46.719 ;
        RECT  1.026 46.161 73.656 46.179 ;
        RECT  1.026 45.621 73.656 45.639 ;
        RECT  1.026 45.081 73.656 45.099 ;
        RECT  1.026 44.541 73.656 44.559 ;
        RECT  1.026 44.001 73.656 44.019 ;
        RECT  1.026 43.461 73.656 43.479 ;
        RECT  1.026 42.921 73.656 42.939 ;
        RECT  1.026 42.381 73.656 42.399 ;
        RECT  1.026 41.841 73.656 41.859 ;
        RECT  1.026 41.301 73.656 41.319 ;
        RECT  1.026 40.761 73.656 40.779 ;
        RECT  1.026 40.221 73.656 40.239 ;
        RECT  1.026 39.681 73.656 39.699 ;
        RECT  1.026 39.141 73.656 39.159 ;
        RECT  1.026 38.601 73.656 38.619 ;
        RECT  1.026 38.061 73.656 38.079 ;
        RECT  1.026 37.521 73.656 37.539 ;
        RECT  1.026 36.981 73.656 36.999 ;
        RECT  1.026 36.441 73.656 36.459 ;
        RECT  1.026 35.901 73.656 35.919 ;
        RECT  1.026 35.361 73.656 35.379 ;
        RECT  1.026 34.821 73.656 34.839 ;
        RECT  1.026 34.281 73.656 34.299 ;
        RECT  1.026 33.741 73.656 33.759 ;
        RECT  1.026 33.201 73.656 33.219 ;
        RECT  1.026 32.661 73.656 32.679 ;
        RECT  1.026 32.121 73.656 32.139 ;
        RECT  1.026 31.581 73.656 31.599 ;
        RECT  1.026 31.041 73.656 31.059 ;
        RECT  1.026 30.501 73.656 30.519 ;
        RECT  1.026 29.961 73.656 29.979 ;
        RECT  1.026 29.421 73.656 29.439 ;
        RECT  1.026 28.881 73.656 28.899 ;
        RECT  1.026 28.341 73.656 28.359 ;
        RECT  1.026 27.801 73.656 27.819 ;
        RECT  1.026 27.261 73.656 27.279 ;
        RECT  1.026 26.721 73.656 26.739 ;
        RECT  1.026 26.181 73.656 26.199 ;
        RECT  1.026 25.641 73.656 25.659 ;
        RECT  1.026 25.101 73.656 25.119 ;
        RECT  1.026 24.561 73.656 24.579 ;
        RECT  1.026 24.021 73.656 24.039 ;
        RECT  1.026 23.481 73.656 23.499 ;
        RECT  1.026 22.941 73.656 22.959 ;
        RECT  1.026 22.401 73.656 22.419 ;
        RECT  1.026 21.861 73.656 21.879 ;
        RECT  1.026 21.321 73.656 21.339 ;
        RECT  1.026 20.781 73.656 20.799 ;
        RECT  1.026 20.241 73.656 20.259 ;
        RECT  1.026 19.701 73.656 19.719 ;
        RECT  1.026 19.161 73.656 19.179 ;
        RECT  1.026 18.621 73.656 18.639 ;
        RECT  1.026 18.081 73.656 18.099 ;
        RECT  1.026 17.541 73.656 17.559 ;
        RECT  1.026 17.001 73.656 17.019 ;
        RECT  1.026 16.461 73.656 16.479 ;
        RECT  1.026 15.921 73.656 15.939 ;
        RECT  1.026 15.381 73.656 15.399 ;
        RECT  1.026 14.841 73.656 14.859 ;
        RECT  1.026 14.301 73.656 14.319 ;
        RECT  1.026 13.761 73.656 13.779 ;
        RECT  1.026 13.221 73.656 13.239 ;
        RECT  1.026 12.681 73.656 12.699 ;
        RECT  1.026 12.141 73.656 12.159 ;
        RECT  1.026 11.601 73.656 11.619 ;
        RECT  1.026 11.061 73.656 11.079 ;
        RECT  1.026 10.521 73.656 10.539 ;
        RECT  1.026 9.981 73.656 9.999 ;
        RECT  1.026 9.441 73.656 9.459 ;
        RECT  1.026 8.901 73.656 8.919 ;
        RECT  1.026 8.361 73.656 8.379 ;
        RECT  1.026 7.821 73.656 7.839 ;
        RECT  1.026 7.281 73.656 7.299 ;
        RECT  1.026 6.741 73.656 6.759 ;
        RECT  1.026 6.201 73.656 6.219 ;
        RECT  1.026 5.661 73.656 5.679 ;
        RECT  1.026 5.121 73.656 5.139 ;
        RECT  1.026 4.581 73.656 4.599 ;
        RECT  1.026 4.041 73.656 4.059 ;
        RECT  1.026 3.501 73.656 3.519 ;
        RECT  1.026 2.961 73.656 2.979 ;
        RECT  1.026 2.421 73.656 2.439 ;
        RECT  1.026 1.881 73.656 1.899 ;
        RECT  1.026 1.341 73.656 1.359 ;
      LAYER M1 ;
        RECT  1.026 73.161 73.656 73.179 ;
        RECT  1.026 72.621 73.656 72.639 ;
        RECT  1.026 72.081 73.656 72.099 ;
        RECT  1.026 71.541 73.656 71.559 ;
        RECT  1.026 71.001 73.656 71.019 ;
        RECT  1.026 70.461 73.656 70.479 ;
        RECT  1.026 69.921 73.656 69.939 ;
        RECT  1.026 69.381 73.656 69.399 ;
        RECT  1.026 68.841 73.656 68.859 ;
        RECT  1.026 68.301 73.656 68.319 ;
        RECT  1.026 67.761 73.656 67.779 ;
        RECT  1.026 67.221 73.656 67.239 ;
        RECT  1.026 66.681 73.656 66.699 ;
        RECT  1.026 66.141 73.656 66.159 ;
        RECT  1.026 65.601 73.656 65.619 ;
        RECT  1.026 65.061 73.656 65.079 ;
        RECT  1.026 64.521 73.656 64.539 ;
        RECT  1.026 63.981 73.656 63.999 ;
        RECT  1.026 63.441 73.656 63.459 ;
        RECT  1.026 62.901 73.656 62.919 ;
        RECT  1.026 62.361 73.656 62.379 ;
        RECT  1.026 61.821 73.656 61.839 ;
        RECT  1.026 61.281 73.656 61.299 ;
        RECT  1.026 60.741 73.656 60.759 ;
        RECT  1.026 60.201 73.656 60.219 ;
        RECT  1.026 59.661 73.656 59.679 ;
        RECT  1.026 59.121 73.656 59.139 ;
        RECT  1.026 58.581 73.656 58.599 ;
        RECT  1.026 58.041 73.656 58.059 ;
        RECT  1.026 57.501 73.656 57.519 ;
        RECT  1.026 56.961 73.656 56.979 ;
        RECT  1.026 56.421 73.656 56.439 ;
        RECT  1.026 55.881 73.656 55.899 ;
        RECT  1.026 55.341 73.656 55.359 ;
        RECT  1.026 54.801 73.656 54.819 ;
        RECT  1.026 54.261 73.656 54.279 ;
        RECT  1.026 53.721 73.656 53.739 ;
        RECT  1.026 53.181 73.656 53.199 ;
        RECT  1.026 52.641 73.656 52.659 ;
        RECT  1.026 52.101 73.656 52.119 ;
        RECT  1.026 51.561 73.656 51.579 ;
        RECT  1.026 51.021 73.656 51.039 ;
        RECT  1.026 50.481 73.656 50.499 ;
        RECT  1.026 49.941 73.656 49.959 ;
        RECT  1.026 49.401 73.656 49.419 ;
        RECT  1.026 48.861 73.656 48.879 ;
        RECT  1.026 48.321 73.656 48.339 ;
        RECT  1.026 47.781 73.656 47.799 ;
        RECT  1.026 47.241 73.656 47.259 ;
        RECT  1.026 46.701 73.656 46.719 ;
        RECT  1.026 46.161 73.656 46.179 ;
        RECT  1.026 45.621 73.656 45.639 ;
        RECT  1.026 45.081 73.656 45.099 ;
        RECT  1.026 44.541 73.656 44.559 ;
        RECT  1.026 44.001 73.656 44.019 ;
        RECT  1.026 43.461 73.656 43.479 ;
        RECT  1.026 42.921 73.656 42.939 ;
        RECT  1.026 42.381 73.656 42.399 ;
        RECT  1.026 41.841 73.656 41.859 ;
        RECT  1.026 41.301 73.656 41.319 ;
        RECT  1.026 40.761 73.656 40.779 ;
        RECT  1.026 40.221 73.656 40.239 ;
        RECT  1.026 39.681 73.656 39.699 ;
        RECT  1.026 39.141 73.656 39.159 ;
        RECT  1.026 38.601 73.656 38.619 ;
        RECT  1.026 38.061 73.656 38.079 ;
        RECT  1.026 37.521 73.656 37.539 ;
        RECT  1.026 36.981 73.656 36.999 ;
        RECT  1.026 36.441 73.656 36.459 ;
        RECT  1.026 35.901 73.656 35.919 ;
        RECT  1.026 35.361 73.656 35.379 ;
        RECT  1.026 34.821 73.656 34.839 ;
        RECT  1.026 34.281 73.656 34.299 ;
        RECT  1.026 33.741 73.656 33.759 ;
        RECT  1.026 33.201 73.656 33.219 ;
        RECT  1.026 32.661 73.656 32.679 ;
        RECT  1.026 32.121 73.656 32.139 ;
        RECT  1.026 31.581 73.656 31.599 ;
        RECT  1.026 31.041 73.656 31.059 ;
        RECT  1.026 30.501 73.656 30.519 ;
        RECT  1.026 29.961 73.656 29.979 ;
        RECT  1.026 29.421 73.656 29.439 ;
        RECT  1.026 28.881 73.656 28.899 ;
        RECT  1.026 28.341 73.656 28.359 ;
        RECT  1.026 27.801 73.656 27.819 ;
        RECT  1.026 27.261 73.656 27.279 ;
        RECT  1.026 26.721 73.656 26.739 ;
        RECT  1.026 26.181 73.656 26.199 ;
        RECT  1.026 25.641 73.656 25.659 ;
        RECT  1.026 25.101 73.656 25.119 ;
        RECT  1.026 24.561 73.656 24.579 ;
        RECT  1.026 24.021 73.656 24.039 ;
        RECT  1.026 23.481 73.656 23.499 ;
        RECT  1.026 22.941 73.656 22.959 ;
        RECT  1.026 22.401 73.656 22.419 ;
        RECT  1.026 21.861 73.656 21.879 ;
        RECT  1.026 21.321 73.656 21.339 ;
        RECT  1.026 20.781 73.656 20.799 ;
        RECT  1.026 20.241 73.656 20.259 ;
        RECT  1.026 19.701 73.656 19.719 ;
        RECT  1.026 19.161 73.656 19.179 ;
        RECT  1.026 18.621 73.656 18.639 ;
        RECT  1.026 18.081 73.656 18.099 ;
        RECT  1.026 17.541 73.656 17.559 ;
        RECT  1.026 17.001 73.656 17.019 ;
        RECT  1.026 16.461 73.656 16.479 ;
        RECT  1.026 15.921 73.656 15.939 ;
        RECT  1.026 15.381 73.656 15.399 ;
        RECT  1.026 14.841 73.656 14.859 ;
        RECT  1.026 14.301 73.656 14.319 ;
        RECT  1.026 13.761 73.656 13.779 ;
        RECT  1.026 13.221 73.656 13.239 ;
        RECT  1.026 12.681 73.656 12.699 ;
        RECT  1.026 12.141 73.656 12.159 ;
        RECT  1.026 11.601 73.656 11.619 ;
        RECT  1.026 11.061 73.656 11.079 ;
        RECT  1.026 10.521 73.656 10.539 ;
        RECT  1.026 9.981 73.656 9.999 ;
        RECT  1.026 9.441 73.656 9.459 ;
        RECT  1.026 8.901 73.656 8.919 ;
        RECT  1.026 8.361 73.656 8.379 ;
        RECT  1.026 7.821 73.656 7.839 ;
        RECT  1.026 7.281 73.656 7.299 ;
        RECT  1.026 6.741 73.656 6.759 ;
        RECT  1.026 6.201 73.656 6.219 ;
        RECT  1.026 5.661 73.656 5.679 ;
        RECT  1.026 5.121 73.656 5.139 ;
        RECT  1.026 4.581 73.656 4.599 ;
        RECT  1.026 4.041 73.656 4.059 ;
        RECT  1.026 3.501 73.656 3.519 ;
        RECT  1.026 2.961 73.656 2.979 ;
        RECT  1.026 2.421 73.656 2.439 ;
        RECT  1.026 1.881 73.656 1.899 ;
        RECT  1.026 1.341 73.656 1.359 ;
      VIA 72.366 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.462 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.558 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 67.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 61.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.366 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 73.153 72.411 73.187 ;
      VIA 72.366 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 72.613 72.411 72.647 ;
      VIA 72.366 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 72.073 72.411 72.107 ;
      VIA 72.366 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 71.533 72.411 71.567 ;
      VIA 72.366 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 70.993 72.411 71.027 ;
      VIA 72.366 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 70.453 72.411 70.487 ;
      VIA 72.366 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 69.913 72.411 69.947 ;
      VIA 72.366 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 69.373 72.411 69.407 ;
      VIA 72.366 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 68.833 72.411 68.867 ;
      VIA 72.366 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 68.293 72.411 68.327 ;
      VIA 72.366 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 67.753 72.411 67.787 ;
      VIA 72.366 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 67.213 72.411 67.247 ;
      VIA 72.366 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 66.673 72.411 66.707 ;
      VIA 72.366 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 66.133 72.411 66.167 ;
      VIA 72.366 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 65.593 72.411 65.627 ;
      VIA 72.366 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 65.053 72.411 65.087 ;
      VIA 72.366 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 64.513 72.411 64.547 ;
      VIA 72.366 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 63.973 72.411 64.007 ;
      VIA 72.366 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 63.433 72.411 63.467 ;
      VIA 72.366 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 62.893 72.411 62.927 ;
      VIA 72.366 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 62.353 72.411 62.387 ;
      VIA 72.366 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 61.813 72.411 61.847 ;
      VIA 72.366 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 61.273 72.411 61.307 ;
      VIA 72.366 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 60.733 72.411 60.767 ;
      VIA 72.366 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 60.193 72.411 60.227 ;
      VIA 72.366 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 59.653 72.411 59.687 ;
      VIA 72.366 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 59.113 72.411 59.147 ;
      VIA 72.366 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 58.573 72.411 58.607 ;
      VIA 72.366 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 58.033 72.411 58.067 ;
      VIA 72.366 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 57.493 72.411 57.527 ;
      VIA 72.366 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 56.953 72.411 56.987 ;
      VIA 72.366 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 56.413 72.411 56.447 ;
      VIA 72.366 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 55.873 72.411 55.907 ;
      VIA 72.366 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 55.333 72.411 55.367 ;
      VIA 72.366 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 54.793 72.411 54.827 ;
      VIA 72.366 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 54.253 72.411 54.287 ;
      VIA 72.366 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 53.713 72.411 53.747 ;
      VIA 72.366 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 53.173 72.411 53.207 ;
      VIA 72.366 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 52.633 72.411 52.667 ;
      VIA 72.366 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 52.093 72.411 52.127 ;
      VIA 72.366 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 51.553 72.411 51.587 ;
      VIA 72.366 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 51.013 72.411 51.047 ;
      VIA 72.366 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 50.473 72.411 50.507 ;
      VIA 72.366 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 49.933 72.411 49.967 ;
      VIA 72.366 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 49.393 72.411 49.427 ;
      VIA 72.366 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 48.853 72.411 48.887 ;
      VIA 72.366 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 48.313 72.411 48.347 ;
      VIA 72.366 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 47.773 72.411 47.807 ;
      VIA 72.366 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 47.233 72.411 47.267 ;
      VIA 72.366 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 46.693 72.411 46.727 ;
      VIA 72.366 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 46.153 72.411 46.187 ;
      VIA 72.366 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 45.613 72.411 45.647 ;
      VIA 72.366 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 45.073 72.411 45.107 ;
      VIA 72.366 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 44.533 72.411 44.567 ;
      VIA 72.366 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 43.993 72.411 44.027 ;
      VIA 72.366 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 43.453 72.411 43.487 ;
      VIA 72.366 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 42.913 72.411 42.947 ;
      VIA 72.366 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 42.373 72.411 42.407 ;
      VIA 72.366 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 41.833 72.411 41.867 ;
      VIA 72.366 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 41.293 72.411 41.327 ;
      VIA 72.366 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 40.753 72.411 40.787 ;
      VIA 72.366 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 40.213 72.411 40.247 ;
      VIA 72.366 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 39.673 72.411 39.707 ;
      VIA 72.366 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 39.133 72.411 39.167 ;
      VIA 72.366 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 38.593 72.411 38.627 ;
      VIA 72.366 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 38.053 72.411 38.087 ;
      VIA 72.366 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 37.513 72.411 37.547 ;
      VIA 72.366 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 36.973 72.411 37.007 ;
      VIA 72.366 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 36.433 72.411 36.467 ;
      VIA 72.366 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 35.893 72.411 35.927 ;
      VIA 72.366 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 35.353 72.411 35.387 ;
      VIA 72.366 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 34.813 72.411 34.847 ;
      VIA 72.366 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 34.273 72.411 34.307 ;
      VIA 72.366 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 33.733 72.411 33.767 ;
      VIA 72.366 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 33.193 72.411 33.227 ;
      VIA 72.366 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 32.653 72.411 32.687 ;
      VIA 72.366 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 32.113 72.411 32.147 ;
      VIA 72.366 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 31.573 72.411 31.607 ;
      VIA 72.366 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 31.033 72.411 31.067 ;
      VIA 72.366 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 30.493 72.411 30.527 ;
      VIA 72.366 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 29.953 72.411 29.987 ;
      VIA 72.366 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 29.413 72.411 29.447 ;
      VIA 72.366 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 28.873 72.411 28.907 ;
      VIA 72.366 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 28.333 72.411 28.367 ;
      VIA 72.366 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 27.793 72.411 27.827 ;
      VIA 72.366 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 27.253 72.411 27.287 ;
      VIA 72.366 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 26.713 72.411 26.747 ;
      VIA 72.366 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 26.173 72.411 26.207 ;
      VIA 72.366 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 25.633 72.411 25.667 ;
      VIA 72.366 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 25.093 72.411 25.127 ;
      VIA 72.366 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 24.553 72.411 24.587 ;
      VIA 72.366 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 24.013 72.411 24.047 ;
      VIA 72.366 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 23.473 72.411 23.507 ;
      VIA 72.366 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 22.933 72.411 22.967 ;
      VIA 72.366 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 22.393 72.411 22.427 ;
      VIA 72.366 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 21.853 72.411 21.887 ;
      VIA 72.366 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 21.313 72.411 21.347 ;
      VIA 72.366 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 20.773 72.411 20.807 ;
      VIA 72.366 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 20.233 72.411 20.267 ;
      VIA 72.366 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 19.693 72.411 19.727 ;
      VIA 72.366 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 19.153 72.411 19.187 ;
      VIA 72.366 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 18.613 72.411 18.647 ;
      VIA 72.366 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 18.073 72.411 18.107 ;
      VIA 72.366 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 17.533 72.411 17.567 ;
      VIA 72.366 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 16.993 72.411 17.027 ;
      VIA 72.366 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 16.453 72.411 16.487 ;
      VIA 72.366 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 15.913 72.411 15.947 ;
      VIA 72.366 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 15.373 72.411 15.407 ;
      VIA 72.366 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 14.833 72.411 14.867 ;
      VIA 72.366 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 14.293 72.411 14.327 ;
      VIA 72.366 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 13.753 72.411 13.787 ;
      VIA 72.366 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 13.213 72.411 13.247 ;
      VIA 72.366 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 12.673 72.411 12.707 ;
      VIA 72.366 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 12.133 72.411 12.167 ;
      VIA 72.366 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 11.593 72.411 11.627 ;
      VIA 72.366 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 11.053 72.411 11.087 ;
      VIA 72.366 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 10.513 72.411 10.547 ;
      VIA 72.366 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 9.973 72.411 10.007 ;
      VIA 72.366 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 9.433 72.411 9.467 ;
      VIA 72.366 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 8.893 72.411 8.927 ;
      VIA 72.366 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 8.353 72.411 8.387 ;
      VIA 72.366 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 7.813 72.411 7.847 ;
      VIA 72.366 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 7.273 72.411 7.307 ;
      VIA 72.366 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 6.733 72.411 6.767 ;
      VIA 72.366 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 6.193 72.411 6.227 ;
      VIA 72.366 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 5.653 72.411 5.687 ;
      VIA 72.366 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 5.113 72.411 5.147 ;
      VIA 72.366 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 4.573 72.411 4.607 ;
      VIA 72.366 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 4.033 72.411 4.067 ;
      VIA 72.366 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 3.493 72.411 3.527 ;
      VIA 72.366 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 2.953 72.411 2.987 ;
      VIA 72.366 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 2.413 72.411 2.447 ;
      VIA 72.366 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 1.873 72.411 1.907 ;
      VIA 72.366 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.366 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.321 1.333 72.411 1.367 ;
      VIA 72.366 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.366 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 73.153 66.507 73.187 ;
      VIA 66.462 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 72.613 66.507 72.647 ;
      VIA 66.462 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 72.073 66.507 72.107 ;
      VIA 66.462 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 71.533 66.507 71.567 ;
      VIA 66.462 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 70.993 66.507 71.027 ;
      VIA 66.462 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 70.453 66.507 70.487 ;
      VIA 66.462 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 69.913 66.507 69.947 ;
      VIA 66.462 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 69.373 66.507 69.407 ;
      VIA 66.462 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 68.833 66.507 68.867 ;
      VIA 66.462 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 68.293 66.507 68.327 ;
      VIA 66.462 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 67.753 66.507 67.787 ;
      VIA 66.462 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 67.213 66.507 67.247 ;
      VIA 66.462 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 66.673 66.507 66.707 ;
      VIA 66.462 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 66.133 66.507 66.167 ;
      VIA 66.462 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 65.593 66.507 65.627 ;
      VIA 66.462 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 65.053 66.507 65.087 ;
      VIA 66.462 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 64.513 66.507 64.547 ;
      VIA 66.462 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 63.973 66.507 64.007 ;
      VIA 66.462 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 63.433 66.507 63.467 ;
      VIA 66.462 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 62.893 66.507 62.927 ;
      VIA 66.462 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 62.353 66.507 62.387 ;
      VIA 66.462 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 61.813 66.507 61.847 ;
      VIA 66.462 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 61.273 66.507 61.307 ;
      VIA 66.462 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 60.733 66.507 60.767 ;
      VIA 66.462 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 60.193 66.507 60.227 ;
      VIA 66.462 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 59.653 66.507 59.687 ;
      VIA 66.462 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 59.113 66.507 59.147 ;
      VIA 66.462 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 58.573 66.507 58.607 ;
      VIA 66.462 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 58.033 66.507 58.067 ;
      VIA 66.462 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 57.493 66.507 57.527 ;
      VIA 66.462 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 56.953 66.507 56.987 ;
      VIA 66.462 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 56.413 66.507 56.447 ;
      VIA 66.462 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 55.873 66.507 55.907 ;
      VIA 66.462 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 55.333 66.507 55.367 ;
      VIA 66.462 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 54.793 66.507 54.827 ;
      VIA 66.462 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 54.253 66.507 54.287 ;
      VIA 66.462 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 53.713 66.507 53.747 ;
      VIA 66.462 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 53.173 66.507 53.207 ;
      VIA 66.462 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 52.633 66.507 52.667 ;
      VIA 66.462 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 52.093 66.507 52.127 ;
      VIA 66.462 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 51.553 66.507 51.587 ;
      VIA 66.462 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 51.013 66.507 51.047 ;
      VIA 66.462 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 50.473 66.507 50.507 ;
      VIA 66.462 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 49.933 66.507 49.967 ;
      VIA 66.462 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 49.393 66.507 49.427 ;
      VIA 66.462 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 48.853 66.507 48.887 ;
      VIA 66.462 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 48.313 66.507 48.347 ;
      VIA 66.462 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 47.773 66.507 47.807 ;
      VIA 66.462 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 47.233 66.507 47.267 ;
      VIA 66.462 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 46.693 66.507 46.727 ;
      VIA 66.462 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 46.153 66.507 46.187 ;
      VIA 66.462 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 45.613 66.507 45.647 ;
      VIA 66.462 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 45.073 66.507 45.107 ;
      VIA 66.462 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 44.533 66.507 44.567 ;
      VIA 66.462 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 43.993 66.507 44.027 ;
      VIA 66.462 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 43.453 66.507 43.487 ;
      VIA 66.462 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 42.913 66.507 42.947 ;
      VIA 66.462 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 42.373 66.507 42.407 ;
      VIA 66.462 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 41.833 66.507 41.867 ;
      VIA 66.462 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 41.293 66.507 41.327 ;
      VIA 66.462 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 40.753 66.507 40.787 ;
      VIA 66.462 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 40.213 66.507 40.247 ;
      VIA 66.462 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 39.673 66.507 39.707 ;
      VIA 66.462 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 39.133 66.507 39.167 ;
      VIA 66.462 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 38.593 66.507 38.627 ;
      VIA 66.462 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 38.053 66.507 38.087 ;
      VIA 66.462 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 37.513 66.507 37.547 ;
      VIA 66.462 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 36.973 66.507 37.007 ;
      VIA 66.462 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 36.433 66.507 36.467 ;
      VIA 66.462 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 35.893 66.507 35.927 ;
      VIA 66.462 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 35.353 66.507 35.387 ;
      VIA 66.462 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 34.813 66.507 34.847 ;
      VIA 66.462 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 34.273 66.507 34.307 ;
      VIA 66.462 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 33.733 66.507 33.767 ;
      VIA 66.462 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 33.193 66.507 33.227 ;
      VIA 66.462 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 32.653 66.507 32.687 ;
      VIA 66.462 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 32.113 66.507 32.147 ;
      VIA 66.462 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 31.573 66.507 31.607 ;
      VIA 66.462 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 31.033 66.507 31.067 ;
      VIA 66.462 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 30.493 66.507 30.527 ;
      VIA 66.462 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 29.953 66.507 29.987 ;
      VIA 66.462 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 29.413 66.507 29.447 ;
      VIA 66.462 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 28.873 66.507 28.907 ;
      VIA 66.462 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 28.333 66.507 28.367 ;
      VIA 66.462 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 27.793 66.507 27.827 ;
      VIA 66.462 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 27.253 66.507 27.287 ;
      VIA 66.462 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 26.713 66.507 26.747 ;
      VIA 66.462 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 26.173 66.507 26.207 ;
      VIA 66.462 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 25.633 66.507 25.667 ;
      VIA 66.462 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 25.093 66.507 25.127 ;
      VIA 66.462 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 24.553 66.507 24.587 ;
      VIA 66.462 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 24.013 66.507 24.047 ;
      VIA 66.462 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 23.473 66.507 23.507 ;
      VIA 66.462 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 22.933 66.507 22.967 ;
      VIA 66.462 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 22.393 66.507 22.427 ;
      VIA 66.462 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 21.853 66.507 21.887 ;
      VIA 66.462 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 21.313 66.507 21.347 ;
      VIA 66.462 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 20.773 66.507 20.807 ;
      VIA 66.462 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 20.233 66.507 20.267 ;
      VIA 66.462 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 19.693 66.507 19.727 ;
      VIA 66.462 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 19.153 66.507 19.187 ;
      VIA 66.462 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 18.613 66.507 18.647 ;
      VIA 66.462 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 18.073 66.507 18.107 ;
      VIA 66.462 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 17.533 66.507 17.567 ;
      VIA 66.462 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 16.993 66.507 17.027 ;
      VIA 66.462 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 16.453 66.507 16.487 ;
      VIA 66.462 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 15.913 66.507 15.947 ;
      VIA 66.462 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 15.373 66.507 15.407 ;
      VIA 66.462 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 14.833 66.507 14.867 ;
      VIA 66.462 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 14.293 66.507 14.327 ;
      VIA 66.462 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 13.753 66.507 13.787 ;
      VIA 66.462 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 13.213 66.507 13.247 ;
      VIA 66.462 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 12.673 66.507 12.707 ;
      VIA 66.462 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 12.133 66.507 12.167 ;
      VIA 66.462 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 11.593 66.507 11.627 ;
      VIA 66.462 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 11.053 66.507 11.087 ;
      VIA 66.462 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 10.513 66.507 10.547 ;
      VIA 66.462 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 9.973 66.507 10.007 ;
      VIA 66.462 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 9.433 66.507 9.467 ;
      VIA 66.462 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 8.893 66.507 8.927 ;
      VIA 66.462 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 8.353 66.507 8.387 ;
      VIA 66.462 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 7.813 66.507 7.847 ;
      VIA 66.462 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 7.273 66.507 7.307 ;
      VIA 66.462 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 6.733 66.507 6.767 ;
      VIA 66.462 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 6.193 66.507 6.227 ;
      VIA 66.462 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 5.653 66.507 5.687 ;
      VIA 66.462 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 5.113 66.507 5.147 ;
      VIA 66.462 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 4.573 66.507 4.607 ;
      VIA 66.462 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 4.033 66.507 4.067 ;
      VIA 66.462 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 3.493 66.507 3.527 ;
      VIA 66.462 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 2.953 66.507 2.987 ;
      VIA 66.462 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 2.413 66.507 2.447 ;
      VIA 66.462 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 1.873 66.507 1.907 ;
      VIA 66.462 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.462 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.417 1.333 66.507 1.367 ;
      VIA 66.462 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.462 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 73.153 60.603 73.187 ;
      VIA 60.558 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 72.613 60.603 72.647 ;
      VIA 60.558 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 72.073 60.603 72.107 ;
      VIA 60.558 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 71.533 60.603 71.567 ;
      VIA 60.558 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 70.993 60.603 71.027 ;
      VIA 60.558 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 70.453 60.603 70.487 ;
      VIA 60.558 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 69.913 60.603 69.947 ;
      VIA 60.558 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 69.373 60.603 69.407 ;
      VIA 60.558 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 68.833 60.603 68.867 ;
      VIA 60.558 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 68.293 60.603 68.327 ;
      VIA 60.558 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 67.753 60.603 67.787 ;
      VIA 60.558 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 67.213 60.603 67.247 ;
      VIA 60.558 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 66.673 60.603 66.707 ;
      VIA 60.558 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 66.133 60.603 66.167 ;
      VIA 60.558 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 65.593 60.603 65.627 ;
      VIA 60.558 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 65.053 60.603 65.087 ;
      VIA 60.558 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 64.513 60.603 64.547 ;
      VIA 60.558 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 63.973 60.603 64.007 ;
      VIA 60.558 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 63.433 60.603 63.467 ;
      VIA 60.558 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 62.893 60.603 62.927 ;
      VIA 60.558 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 62.353 60.603 62.387 ;
      VIA 60.558 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 61.813 60.603 61.847 ;
      VIA 60.558 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 61.273 60.603 61.307 ;
      VIA 60.558 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 60.733 60.603 60.767 ;
      VIA 60.558 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 60.193 60.603 60.227 ;
      VIA 60.558 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 59.653 60.603 59.687 ;
      VIA 60.558 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 59.113 60.603 59.147 ;
      VIA 60.558 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 58.573 60.603 58.607 ;
      VIA 60.558 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 58.033 60.603 58.067 ;
      VIA 60.558 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 57.493 60.603 57.527 ;
      VIA 60.558 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 56.953 60.603 56.987 ;
      VIA 60.558 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 56.413 60.603 56.447 ;
      VIA 60.558 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 55.873 60.603 55.907 ;
      VIA 60.558 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 55.333 60.603 55.367 ;
      VIA 60.558 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 54.793 60.603 54.827 ;
      VIA 60.558 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 54.253 60.603 54.287 ;
      VIA 60.558 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 53.713 60.603 53.747 ;
      VIA 60.558 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 53.173 60.603 53.207 ;
      VIA 60.558 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 52.633 60.603 52.667 ;
      VIA 60.558 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 52.093 60.603 52.127 ;
      VIA 60.558 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 51.553 60.603 51.587 ;
      VIA 60.558 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 51.013 60.603 51.047 ;
      VIA 60.558 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 50.473 60.603 50.507 ;
      VIA 60.558 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 49.933 60.603 49.967 ;
      VIA 60.558 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 49.393 60.603 49.427 ;
      VIA 60.558 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 48.853 60.603 48.887 ;
      VIA 60.558 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 48.313 60.603 48.347 ;
      VIA 60.558 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 47.773 60.603 47.807 ;
      VIA 60.558 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 47.233 60.603 47.267 ;
      VIA 60.558 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 46.693 60.603 46.727 ;
      VIA 60.558 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 46.153 60.603 46.187 ;
      VIA 60.558 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 45.613 60.603 45.647 ;
      VIA 60.558 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 45.073 60.603 45.107 ;
      VIA 60.558 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 44.533 60.603 44.567 ;
      VIA 60.558 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 43.993 60.603 44.027 ;
      VIA 60.558 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 43.453 60.603 43.487 ;
      VIA 60.558 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 42.913 60.603 42.947 ;
      VIA 60.558 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 42.373 60.603 42.407 ;
      VIA 60.558 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 41.833 60.603 41.867 ;
      VIA 60.558 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 41.293 60.603 41.327 ;
      VIA 60.558 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 40.753 60.603 40.787 ;
      VIA 60.558 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 40.213 60.603 40.247 ;
      VIA 60.558 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 39.673 60.603 39.707 ;
      VIA 60.558 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 39.133 60.603 39.167 ;
      VIA 60.558 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 38.593 60.603 38.627 ;
      VIA 60.558 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 38.053 60.603 38.087 ;
      VIA 60.558 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 37.513 60.603 37.547 ;
      VIA 60.558 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 36.973 60.603 37.007 ;
      VIA 60.558 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 36.433 60.603 36.467 ;
      VIA 60.558 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 35.893 60.603 35.927 ;
      VIA 60.558 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 35.353 60.603 35.387 ;
      VIA 60.558 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 34.813 60.603 34.847 ;
      VIA 60.558 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 34.273 60.603 34.307 ;
      VIA 60.558 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 33.733 60.603 33.767 ;
      VIA 60.558 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 33.193 60.603 33.227 ;
      VIA 60.558 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 32.653 60.603 32.687 ;
      VIA 60.558 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 32.113 60.603 32.147 ;
      VIA 60.558 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 31.573 60.603 31.607 ;
      VIA 60.558 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 31.033 60.603 31.067 ;
      VIA 60.558 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 30.493 60.603 30.527 ;
      VIA 60.558 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 29.953 60.603 29.987 ;
      VIA 60.558 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 29.413 60.603 29.447 ;
      VIA 60.558 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 28.873 60.603 28.907 ;
      VIA 60.558 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 28.333 60.603 28.367 ;
      VIA 60.558 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 27.793 60.603 27.827 ;
      VIA 60.558 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 27.253 60.603 27.287 ;
      VIA 60.558 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 26.713 60.603 26.747 ;
      VIA 60.558 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 26.173 60.603 26.207 ;
      VIA 60.558 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 25.633 60.603 25.667 ;
      VIA 60.558 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 25.093 60.603 25.127 ;
      VIA 60.558 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 24.553 60.603 24.587 ;
      VIA 60.558 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 24.013 60.603 24.047 ;
      VIA 60.558 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 23.473 60.603 23.507 ;
      VIA 60.558 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 22.933 60.603 22.967 ;
      VIA 60.558 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 22.393 60.603 22.427 ;
      VIA 60.558 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 21.853 60.603 21.887 ;
      VIA 60.558 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 21.313 60.603 21.347 ;
      VIA 60.558 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 20.773 60.603 20.807 ;
      VIA 60.558 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 20.233 60.603 20.267 ;
      VIA 60.558 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 19.693 60.603 19.727 ;
      VIA 60.558 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 19.153 60.603 19.187 ;
      VIA 60.558 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 18.613 60.603 18.647 ;
      VIA 60.558 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 18.073 60.603 18.107 ;
      VIA 60.558 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 17.533 60.603 17.567 ;
      VIA 60.558 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 16.993 60.603 17.027 ;
      VIA 60.558 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 16.453 60.603 16.487 ;
      VIA 60.558 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 15.913 60.603 15.947 ;
      VIA 60.558 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 15.373 60.603 15.407 ;
      VIA 60.558 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 14.833 60.603 14.867 ;
      VIA 60.558 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 14.293 60.603 14.327 ;
      VIA 60.558 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 13.753 60.603 13.787 ;
      VIA 60.558 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 13.213 60.603 13.247 ;
      VIA 60.558 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 12.673 60.603 12.707 ;
      VIA 60.558 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 12.133 60.603 12.167 ;
      VIA 60.558 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 11.593 60.603 11.627 ;
      VIA 60.558 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 11.053 60.603 11.087 ;
      VIA 60.558 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 10.513 60.603 10.547 ;
      VIA 60.558 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 9.973 60.603 10.007 ;
      VIA 60.558 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 9.433 60.603 9.467 ;
      VIA 60.558 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 8.893 60.603 8.927 ;
      VIA 60.558 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 8.353 60.603 8.387 ;
      VIA 60.558 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 7.813 60.603 7.847 ;
      VIA 60.558 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 7.273 60.603 7.307 ;
      VIA 60.558 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 6.733 60.603 6.767 ;
      VIA 60.558 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 6.193 60.603 6.227 ;
      VIA 60.558 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 5.653 60.603 5.687 ;
      VIA 60.558 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 5.113 60.603 5.147 ;
      VIA 60.558 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 4.573 60.603 4.607 ;
      VIA 60.558 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 4.033 60.603 4.067 ;
      VIA 60.558 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 3.493 60.603 3.527 ;
      VIA 60.558 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 2.953 60.603 2.987 ;
      VIA 60.558 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 2.413 60.603 2.447 ;
      VIA 60.558 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 1.873 60.603 1.907 ;
      VIA 60.558 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.558 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.513 1.333 60.603 1.367 ;
      VIA 60.558 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.558 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 73.153 54.699 73.187 ;
      VIA 54.654 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 72.613 54.699 72.647 ;
      VIA 54.654 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 72.073 54.699 72.107 ;
      VIA 54.654 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 71.533 54.699 71.567 ;
      VIA 54.654 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 70.993 54.699 71.027 ;
      VIA 54.654 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 70.453 54.699 70.487 ;
      VIA 54.654 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 69.913 54.699 69.947 ;
      VIA 54.654 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 69.373 54.699 69.407 ;
      VIA 54.654 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 68.833 54.699 68.867 ;
      VIA 54.654 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 68.293 54.699 68.327 ;
      VIA 54.654 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 67.753 54.699 67.787 ;
      VIA 54.654 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 67.213 54.699 67.247 ;
      VIA 54.654 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 66.673 54.699 66.707 ;
      VIA 54.654 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 66.133 54.699 66.167 ;
      VIA 54.654 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 65.593 54.699 65.627 ;
      VIA 54.654 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 65.053 54.699 65.087 ;
      VIA 54.654 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 64.513 54.699 64.547 ;
      VIA 54.654 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 63.973 54.699 64.007 ;
      VIA 54.654 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 63.433 54.699 63.467 ;
      VIA 54.654 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 62.893 54.699 62.927 ;
      VIA 54.654 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 62.353 54.699 62.387 ;
      VIA 54.654 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 61.813 54.699 61.847 ;
      VIA 54.654 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 61.273 54.699 61.307 ;
      VIA 54.654 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 60.733 54.699 60.767 ;
      VIA 54.654 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 60.193 54.699 60.227 ;
      VIA 54.654 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 59.653 54.699 59.687 ;
      VIA 54.654 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 59.113 54.699 59.147 ;
      VIA 54.654 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 58.573 54.699 58.607 ;
      VIA 54.654 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 58.033 54.699 58.067 ;
      VIA 54.654 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 57.493 54.699 57.527 ;
      VIA 54.654 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 56.953 54.699 56.987 ;
      VIA 54.654 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 56.413 54.699 56.447 ;
      VIA 54.654 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 55.873 54.699 55.907 ;
      VIA 54.654 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 55.333 54.699 55.367 ;
      VIA 54.654 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 54.793 54.699 54.827 ;
      VIA 54.654 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 54.253 54.699 54.287 ;
      VIA 54.654 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 53.713 54.699 53.747 ;
      VIA 54.654 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 53.173 54.699 53.207 ;
      VIA 54.654 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 52.633 54.699 52.667 ;
      VIA 54.654 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 52.093 54.699 52.127 ;
      VIA 54.654 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 51.553 54.699 51.587 ;
      VIA 54.654 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 51.013 54.699 51.047 ;
      VIA 54.654 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 50.473 54.699 50.507 ;
      VIA 54.654 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 49.933 54.699 49.967 ;
      VIA 54.654 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 49.393 54.699 49.427 ;
      VIA 54.654 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 48.853 54.699 48.887 ;
      VIA 54.654 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 48.313 54.699 48.347 ;
      VIA 54.654 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 47.773 54.699 47.807 ;
      VIA 54.654 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 47.233 54.699 47.267 ;
      VIA 54.654 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 46.693 54.699 46.727 ;
      VIA 54.654 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 46.153 54.699 46.187 ;
      VIA 54.654 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 45.613 54.699 45.647 ;
      VIA 54.654 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 45.073 54.699 45.107 ;
      VIA 54.654 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 44.533 54.699 44.567 ;
      VIA 54.654 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 43.993 54.699 44.027 ;
      VIA 54.654 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 43.453 54.699 43.487 ;
      VIA 54.654 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 42.913 54.699 42.947 ;
      VIA 54.654 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 42.373 54.699 42.407 ;
      VIA 54.654 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 41.833 54.699 41.867 ;
      VIA 54.654 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 41.293 54.699 41.327 ;
      VIA 54.654 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 40.753 54.699 40.787 ;
      VIA 54.654 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 40.213 54.699 40.247 ;
      VIA 54.654 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 39.673 54.699 39.707 ;
      VIA 54.654 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 39.133 54.699 39.167 ;
      VIA 54.654 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 38.593 54.699 38.627 ;
      VIA 54.654 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 38.053 54.699 38.087 ;
      VIA 54.654 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 37.513 54.699 37.547 ;
      VIA 54.654 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 36.973 54.699 37.007 ;
      VIA 54.654 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 36.433 54.699 36.467 ;
      VIA 54.654 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 35.893 54.699 35.927 ;
      VIA 54.654 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 35.353 54.699 35.387 ;
      VIA 54.654 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 34.813 54.699 34.847 ;
      VIA 54.654 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 34.273 54.699 34.307 ;
      VIA 54.654 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 33.733 54.699 33.767 ;
      VIA 54.654 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 33.193 54.699 33.227 ;
      VIA 54.654 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 32.653 54.699 32.687 ;
      VIA 54.654 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 32.113 54.699 32.147 ;
      VIA 54.654 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 31.573 54.699 31.607 ;
      VIA 54.654 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 31.033 54.699 31.067 ;
      VIA 54.654 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 30.493 54.699 30.527 ;
      VIA 54.654 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 29.953 54.699 29.987 ;
      VIA 54.654 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 29.413 54.699 29.447 ;
      VIA 54.654 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 28.873 54.699 28.907 ;
      VIA 54.654 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 28.333 54.699 28.367 ;
      VIA 54.654 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 27.793 54.699 27.827 ;
      VIA 54.654 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 27.253 54.699 27.287 ;
      VIA 54.654 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 26.713 54.699 26.747 ;
      VIA 54.654 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 26.173 54.699 26.207 ;
      VIA 54.654 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 25.633 54.699 25.667 ;
      VIA 54.654 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 25.093 54.699 25.127 ;
      VIA 54.654 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 24.553 54.699 24.587 ;
      VIA 54.654 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 24.013 54.699 24.047 ;
      VIA 54.654 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 23.473 54.699 23.507 ;
      VIA 54.654 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 22.933 54.699 22.967 ;
      VIA 54.654 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 22.393 54.699 22.427 ;
      VIA 54.654 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 21.853 54.699 21.887 ;
      VIA 54.654 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 21.313 54.699 21.347 ;
      VIA 54.654 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 20.773 54.699 20.807 ;
      VIA 54.654 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 20.233 54.699 20.267 ;
      VIA 54.654 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 19.693 54.699 19.727 ;
      VIA 54.654 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 19.153 54.699 19.187 ;
      VIA 54.654 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 18.613 54.699 18.647 ;
      VIA 54.654 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 18.073 54.699 18.107 ;
      VIA 54.654 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 17.533 54.699 17.567 ;
      VIA 54.654 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 16.993 54.699 17.027 ;
      VIA 54.654 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 16.453 54.699 16.487 ;
      VIA 54.654 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 15.913 54.699 15.947 ;
      VIA 54.654 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 15.373 54.699 15.407 ;
      VIA 54.654 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 14.833 54.699 14.867 ;
      VIA 54.654 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 14.293 54.699 14.327 ;
      VIA 54.654 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 13.753 54.699 13.787 ;
      VIA 54.654 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 13.213 54.699 13.247 ;
      VIA 54.654 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 12.673 54.699 12.707 ;
      VIA 54.654 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 12.133 54.699 12.167 ;
      VIA 54.654 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 11.593 54.699 11.627 ;
      VIA 54.654 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 11.053 54.699 11.087 ;
      VIA 54.654 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 10.513 54.699 10.547 ;
      VIA 54.654 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 9.973 54.699 10.007 ;
      VIA 54.654 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 9.433 54.699 9.467 ;
      VIA 54.654 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 8.893 54.699 8.927 ;
      VIA 54.654 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 8.353 54.699 8.387 ;
      VIA 54.654 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 7.813 54.699 7.847 ;
      VIA 54.654 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 7.273 54.699 7.307 ;
      VIA 54.654 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 6.733 54.699 6.767 ;
      VIA 54.654 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 6.193 54.699 6.227 ;
      VIA 54.654 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 5.653 54.699 5.687 ;
      VIA 54.654 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 5.113 54.699 5.147 ;
      VIA 54.654 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 4.573 54.699 4.607 ;
      VIA 54.654 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 4.033 54.699 4.067 ;
      VIA 54.654 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 3.493 54.699 3.527 ;
      VIA 54.654 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 2.953 54.699 2.987 ;
      VIA 54.654 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 2.413 54.699 2.447 ;
      VIA 54.654 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 1.873 54.699 1.907 ;
      VIA 54.654 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 1.333 54.699 1.367 ;
      VIA 54.654 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 73.153 48.795 73.187 ;
      VIA 48.75 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 72.613 48.795 72.647 ;
      VIA 48.75 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 72.073 48.795 72.107 ;
      VIA 48.75 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 71.533 48.795 71.567 ;
      VIA 48.75 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 70.993 48.795 71.027 ;
      VIA 48.75 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 70.453 48.795 70.487 ;
      VIA 48.75 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 69.913 48.795 69.947 ;
      VIA 48.75 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 69.373 48.795 69.407 ;
      VIA 48.75 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 68.833 48.795 68.867 ;
      VIA 48.75 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 68.293 48.795 68.327 ;
      VIA 48.75 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 67.753 48.795 67.787 ;
      VIA 48.75 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 67.213 48.795 67.247 ;
      VIA 48.75 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 66.673 48.795 66.707 ;
      VIA 48.75 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 66.133 48.795 66.167 ;
      VIA 48.75 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 65.593 48.795 65.627 ;
      VIA 48.75 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 65.053 48.795 65.087 ;
      VIA 48.75 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 64.513 48.795 64.547 ;
      VIA 48.75 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 63.973 48.795 64.007 ;
      VIA 48.75 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 63.433 48.795 63.467 ;
      VIA 48.75 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 62.893 48.795 62.927 ;
      VIA 48.75 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 62.353 48.795 62.387 ;
      VIA 48.75 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 61.813 48.795 61.847 ;
      VIA 48.75 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 61.273 48.795 61.307 ;
      VIA 48.75 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 60.733 48.795 60.767 ;
      VIA 48.75 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 60.193 48.795 60.227 ;
      VIA 48.75 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 59.653 48.795 59.687 ;
      VIA 48.75 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 59.113 48.795 59.147 ;
      VIA 48.75 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 58.573 48.795 58.607 ;
      VIA 48.75 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 58.033 48.795 58.067 ;
      VIA 48.75 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 57.493 48.795 57.527 ;
      VIA 48.75 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 56.953 48.795 56.987 ;
      VIA 48.75 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 56.413 48.795 56.447 ;
      VIA 48.75 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 55.873 48.795 55.907 ;
      VIA 48.75 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 55.333 48.795 55.367 ;
      VIA 48.75 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 54.793 48.795 54.827 ;
      VIA 48.75 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 54.253 48.795 54.287 ;
      VIA 48.75 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 53.713 48.795 53.747 ;
      VIA 48.75 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 53.173 48.795 53.207 ;
      VIA 48.75 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 52.633 48.795 52.667 ;
      VIA 48.75 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 52.093 48.795 52.127 ;
      VIA 48.75 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 51.553 48.795 51.587 ;
      VIA 48.75 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 51.013 48.795 51.047 ;
      VIA 48.75 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 50.473 48.795 50.507 ;
      VIA 48.75 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 49.933 48.795 49.967 ;
      VIA 48.75 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 49.393 48.795 49.427 ;
      VIA 48.75 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 48.853 48.795 48.887 ;
      VIA 48.75 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 48.313 48.795 48.347 ;
      VIA 48.75 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 47.773 48.795 47.807 ;
      VIA 48.75 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 47.233 48.795 47.267 ;
      VIA 48.75 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 46.693 48.795 46.727 ;
      VIA 48.75 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 46.153 48.795 46.187 ;
      VIA 48.75 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 45.613 48.795 45.647 ;
      VIA 48.75 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 45.073 48.795 45.107 ;
      VIA 48.75 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 44.533 48.795 44.567 ;
      VIA 48.75 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 43.993 48.795 44.027 ;
      VIA 48.75 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 43.453 48.795 43.487 ;
      VIA 48.75 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 42.913 48.795 42.947 ;
      VIA 48.75 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 42.373 48.795 42.407 ;
      VIA 48.75 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 41.833 48.795 41.867 ;
      VIA 48.75 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 41.293 48.795 41.327 ;
      VIA 48.75 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 40.753 48.795 40.787 ;
      VIA 48.75 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 40.213 48.795 40.247 ;
      VIA 48.75 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 39.673 48.795 39.707 ;
      VIA 48.75 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 39.133 48.795 39.167 ;
      VIA 48.75 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 38.593 48.795 38.627 ;
      VIA 48.75 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 38.053 48.795 38.087 ;
      VIA 48.75 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 37.513 48.795 37.547 ;
      VIA 48.75 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 36.973 48.795 37.007 ;
      VIA 48.75 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 36.433 48.795 36.467 ;
      VIA 48.75 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 35.893 48.795 35.927 ;
      VIA 48.75 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 35.353 48.795 35.387 ;
      VIA 48.75 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 34.813 48.795 34.847 ;
      VIA 48.75 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 34.273 48.795 34.307 ;
      VIA 48.75 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 33.733 48.795 33.767 ;
      VIA 48.75 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 33.193 48.795 33.227 ;
      VIA 48.75 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 32.653 48.795 32.687 ;
      VIA 48.75 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 32.113 48.795 32.147 ;
      VIA 48.75 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 31.573 48.795 31.607 ;
      VIA 48.75 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 31.033 48.795 31.067 ;
      VIA 48.75 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 30.493 48.795 30.527 ;
      VIA 48.75 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 29.953 48.795 29.987 ;
      VIA 48.75 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 29.413 48.795 29.447 ;
      VIA 48.75 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 28.873 48.795 28.907 ;
      VIA 48.75 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 28.333 48.795 28.367 ;
      VIA 48.75 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 27.793 48.795 27.827 ;
      VIA 48.75 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 27.253 48.795 27.287 ;
      VIA 48.75 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 26.713 48.795 26.747 ;
      VIA 48.75 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 26.173 48.795 26.207 ;
      VIA 48.75 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 25.633 48.795 25.667 ;
      VIA 48.75 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 25.093 48.795 25.127 ;
      VIA 48.75 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 24.553 48.795 24.587 ;
      VIA 48.75 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 24.013 48.795 24.047 ;
      VIA 48.75 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 23.473 48.795 23.507 ;
      VIA 48.75 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 22.933 48.795 22.967 ;
      VIA 48.75 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 22.393 48.795 22.427 ;
      VIA 48.75 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 21.853 48.795 21.887 ;
      VIA 48.75 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 21.313 48.795 21.347 ;
      VIA 48.75 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 20.773 48.795 20.807 ;
      VIA 48.75 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 20.233 48.795 20.267 ;
      VIA 48.75 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 19.693 48.795 19.727 ;
      VIA 48.75 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 19.153 48.795 19.187 ;
      VIA 48.75 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 18.613 48.795 18.647 ;
      VIA 48.75 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 18.073 48.795 18.107 ;
      VIA 48.75 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 17.533 48.795 17.567 ;
      VIA 48.75 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 16.993 48.795 17.027 ;
      VIA 48.75 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 16.453 48.795 16.487 ;
      VIA 48.75 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 15.913 48.795 15.947 ;
      VIA 48.75 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 15.373 48.795 15.407 ;
      VIA 48.75 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 14.833 48.795 14.867 ;
      VIA 48.75 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 14.293 48.795 14.327 ;
      VIA 48.75 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 13.753 48.795 13.787 ;
      VIA 48.75 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 13.213 48.795 13.247 ;
      VIA 48.75 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 12.673 48.795 12.707 ;
      VIA 48.75 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 12.133 48.795 12.167 ;
      VIA 48.75 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 11.593 48.795 11.627 ;
      VIA 48.75 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 11.053 48.795 11.087 ;
      VIA 48.75 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 10.513 48.795 10.547 ;
      VIA 48.75 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 9.973 48.795 10.007 ;
      VIA 48.75 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 9.433 48.795 9.467 ;
      VIA 48.75 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 8.893 48.795 8.927 ;
      VIA 48.75 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 8.353 48.795 8.387 ;
      VIA 48.75 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 7.813 48.795 7.847 ;
      VIA 48.75 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 7.273 48.795 7.307 ;
      VIA 48.75 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 6.733 48.795 6.767 ;
      VIA 48.75 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 6.193 48.795 6.227 ;
      VIA 48.75 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 5.653 48.795 5.687 ;
      VIA 48.75 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 5.113 48.795 5.147 ;
      VIA 48.75 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 4.573 48.795 4.607 ;
      VIA 48.75 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 4.033 48.795 4.067 ;
      VIA 48.75 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 3.493 48.795 3.527 ;
      VIA 48.75 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 2.953 48.795 2.987 ;
      VIA 48.75 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 2.413 48.795 2.447 ;
      VIA 48.75 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 1.873 48.795 1.907 ;
      VIA 48.75 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 1.333 48.795 1.367 ;
      VIA 48.75 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 73.153 42.891 73.187 ;
      VIA 42.846 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 72.613 42.891 72.647 ;
      VIA 42.846 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 72.073 42.891 72.107 ;
      VIA 42.846 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 71.533 42.891 71.567 ;
      VIA 42.846 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 70.993 42.891 71.027 ;
      VIA 42.846 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 70.453 42.891 70.487 ;
      VIA 42.846 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 69.913 42.891 69.947 ;
      VIA 42.846 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 69.373 42.891 69.407 ;
      VIA 42.846 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 68.833 42.891 68.867 ;
      VIA 42.846 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 68.293 42.891 68.327 ;
      VIA 42.846 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 67.753 42.891 67.787 ;
      VIA 42.846 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 67.213 42.891 67.247 ;
      VIA 42.846 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 66.673 42.891 66.707 ;
      VIA 42.846 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 66.133 42.891 66.167 ;
      VIA 42.846 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 65.593 42.891 65.627 ;
      VIA 42.846 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 65.053 42.891 65.087 ;
      VIA 42.846 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 64.513 42.891 64.547 ;
      VIA 42.846 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 63.973 42.891 64.007 ;
      VIA 42.846 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 63.433 42.891 63.467 ;
      VIA 42.846 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 62.893 42.891 62.927 ;
      VIA 42.846 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 62.353 42.891 62.387 ;
      VIA 42.846 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 61.813 42.891 61.847 ;
      VIA 42.846 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 61.273 42.891 61.307 ;
      VIA 42.846 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 60.733 42.891 60.767 ;
      VIA 42.846 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 60.193 42.891 60.227 ;
      VIA 42.846 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 59.653 42.891 59.687 ;
      VIA 42.846 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 59.113 42.891 59.147 ;
      VIA 42.846 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 58.573 42.891 58.607 ;
      VIA 42.846 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 58.033 42.891 58.067 ;
      VIA 42.846 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 57.493 42.891 57.527 ;
      VIA 42.846 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 56.953 42.891 56.987 ;
      VIA 42.846 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 56.413 42.891 56.447 ;
      VIA 42.846 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 55.873 42.891 55.907 ;
      VIA 42.846 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 55.333 42.891 55.367 ;
      VIA 42.846 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 54.793 42.891 54.827 ;
      VIA 42.846 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 54.253 42.891 54.287 ;
      VIA 42.846 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 53.713 42.891 53.747 ;
      VIA 42.846 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 53.173 42.891 53.207 ;
      VIA 42.846 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 52.633 42.891 52.667 ;
      VIA 42.846 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 52.093 42.891 52.127 ;
      VIA 42.846 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 51.553 42.891 51.587 ;
      VIA 42.846 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 51.013 42.891 51.047 ;
      VIA 42.846 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 50.473 42.891 50.507 ;
      VIA 42.846 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 49.933 42.891 49.967 ;
      VIA 42.846 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 49.393 42.891 49.427 ;
      VIA 42.846 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 48.853 42.891 48.887 ;
      VIA 42.846 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 48.313 42.891 48.347 ;
      VIA 42.846 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 47.773 42.891 47.807 ;
      VIA 42.846 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 47.233 42.891 47.267 ;
      VIA 42.846 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 46.693 42.891 46.727 ;
      VIA 42.846 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 46.153 42.891 46.187 ;
      VIA 42.846 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 45.613 42.891 45.647 ;
      VIA 42.846 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 45.073 42.891 45.107 ;
      VIA 42.846 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 44.533 42.891 44.567 ;
      VIA 42.846 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 43.993 42.891 44.027 ;
      VIA 42.846 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 43.453 42.891 43.487 ;
      VIA 42.846 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 42.913 42.891 42.947 ;
      VIA 42.846 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 42.373 42.891 42.407 ;
      VIA 42.846 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 41.833 42.891 41.867 ;
      VIA 42.846 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 41.293 42.891 41.327 ;
      VIA 42.846 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 40.753 42.891 40.787 ;
      VIA 42.846 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 40.213 42.891 40.247 ;
      VIA 42.846 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 39.673 42.891 39.707 ;
      VIA 42.846 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 39.133 42.891 39.167 ;
      VIA 42.846 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 38.593 42.891 38.627 ;
      VIA 42.846 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 38.053 42.891 38.087 ;
      VIA 42.846 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 37.513 42.891 37.547 ;
      VIA 42.846 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 36.973 42.891 37.007 ;
      VIA 42.846 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 36.433 42.891 36.467 ;
      VIA 42.846 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 35.893 42.891 35.927 ;
      VIA 42.846 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 35.353 42.891 35.387 ;
      VIA 42.846 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 34.813 42.891 34.847 ;
      VIA 42.846 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 34.273 42.891 34.307 ;
      VIA 42.846 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 33.733 42.891 33.767 ;
      VIA 42.846 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 33.193 42.891 33.227 ;
      VIA 42.846 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 32.653 42.891 32.687 ;
      VIA 42.846 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 32.113 42.891 32.147 ;
      VIA 42.846 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 31.573 42.891 31.607 ;
      VIA 42.846 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 31.033 42.891 31.067 ;
      VIA 42.846 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 30.493 42.891 30.527 ;
      VIA 42.846 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 29.953 42.891 29.987 ;
      VIA 42.846 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 29.413 42.891 29.447 ;
      VIA 42.846 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 28.873 42.891 28.907 ;
      VIA 42.846 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 28.333 42.891 28.367 ;
      VIA 42.846 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 27.793 42.891 27.827 ;
      VIA 42.846 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 27.253 42.891 27.287 ;
      VIA 42.846 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 26.713 42.891 26.747 ;
      VIA 42.846 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 26.173 42.891 26.207 ;
      VIA 42.846 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 25.633 42.891 25.667 ;
      VIA 42.846 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 25.093 42.891 25.127 ;
      VIA 42.846 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 24.553 42.891 24.587 ;
      VIA 42.846 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 24.013 42.891 24.047 ;
      VIA 42.846 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 23.473 42.891 23.507 ;
      VIA 42.846 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 22.933 42.891 22.967 ;
      VIA 42.846 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 22.393 42.891 22.427 ;
      VIA 42.846 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 21.853 42.891 21.887 ;
      VIA 42.846 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 21.313 42.891 21.347 ;
      VIA 42.846 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 20.773 42.891 20.807 ;
      VIA 42.846 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 20.233 42.891 20.267 ;
      VIA 42.846 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 19.693 42.891 19.727 ;
      VIA 42.846 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 19.153 42.891 19.187 ;
      VIA 42.846 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 18.613 42.891 18.647 ;
      VIA 42.846 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 18.073 42.891 18.107 ;
      VIA 42.846 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 17.533 42.891 17.567 ;
      VIA 42.846 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 16.993 42.891 17.027 ;
      VIA 42.846 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 16.453 42.891 16.487 ;
      VIA 42.846 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 15.913 42.891 15.947 ;
      VIA 42.846 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 15.373 42.891 15.407 ;
      VIA 42.846 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 14.833 42.891 14.867 ;
      VIA 42.846 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 14.293 42.891 14.327 ;
      VIA 42.846 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 13.753 42.891 13.787 ;
      VIA 42.846 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 13.213 42.891 13.247 ;
      VIA 42.846 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 12.673 42.891 12.707 ;
      VIA 42.846 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 12.133 42.891 12.167 ;
      VIA 42.846 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 11.593 42.891 11.627 ;
      VIA 42.846 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 11.053 42.891 11.087 ;
      VIA 42.846 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 10.513 42.891 10.547 ;
      VIA 42.846 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 9.973 42.891 10.007 ;
      VIA 42.846 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 9.433 42.891 9.467 ;
      VIA 42.846 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 8.893 42.891 8.927 ;
      VIA 42.846 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 8.353 42.891 8.387 ;
      VIA 42.846 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 7.813 42.891 7.847 ;
      VIA 42.846 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 7.273 42.891 7.307 ;
      VIA 42.846 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 6.733 42.891 6.767 ;
      VIA 42.846 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 6.193 42.891 6.227 ;
      VIA 42.846 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 5.653 42.891 5.687 ;
      VIA 42.846 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 5.113 42.891 5.147 ;
      VIA 42.846 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 4.573 42.891 4.607 ;
      VIA 42.846 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 4.033 42.891 4.067 ;
      VIA 42.846 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 3.493 42.891 3.527 ;
      VIA 42.846 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 2.953 42.891 2.987 ;
      VIA 42.846 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 2.413 42.891 2.447 ;
      VIA 42.846 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 1.873 42.891 1.907 ;
      VIA 42.846 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 1.333 42.891 1.367 ;
      VIA 42.846 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 73.153 36.987 73.187 ;
      VIA 36.942 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 72.613 36.987 72.647 ;
      VIA 36.942 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 72.073 36.987 72.107 ;
      VIA 36.942 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 71.533 36.987 71.567 ;
      VIA 36.942 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 70.993 36.987 71.027 ;
      VIA 36.942 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 70.453 36.987 70.487 ;
      VIA 36.942 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 69.913 36.987 69.947 ;
      VIA 36.942 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 69.373 36.987 69.407 ;
      VIA 36.942 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 68.833 36.987 68.867 ;
      VIA 36.942 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 68.293 36.987 68.327 ;
      VIA 36.942 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 67.753 36.987 67.787 ;
      VIA 36.942 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 67.213 36.987 67.247 ;
      VIA 36.942 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 66.673 36.987 66.707 ;
      VIA 36.942 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 66.133 36.987 66.167 ;
      VIA 36.942 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 65.593 36.987 65.627 ;
      VIA 36.942 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 65.053 36.987 65.087 ;
      VIA 36.942 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 64.513 36.987 64.547 ;
      VIA 36.942 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 63.973 36.987 64.007 ;
      VIA 36.942 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 63.433 36.987 63.467 ;
      VIA 36.942 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 62.893 36.987 62.927 ;
      VIA 36.942 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 62.353 36.987 62.387 ;
      VIA 36.942 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 61.813 36.987 61.847 ;
      VIA 36.942 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 61.273 36.987 61.307 ;
      VIA 36.942 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 60.733 36.987 60.767 ;
      VIA 36.942 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 60.193 36.987 60.227 ;
      VIA 36.942 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 59.653 36.987 59.687 ;
      VIA 36.942 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 59.113 36.987 59.147 ;
      VIA 36.942 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 58.573 36.987 58.607 ;
      VIA 36.942 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 58.033 36.987 58.067 ;
      VIA 36.942 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 57.493 36.987 57.527 ;
      VIA 36.942 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 56.953 36.987 56.987 ;
      VIA 36.942 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 56.413 36.987 56.447 ;
      VIA 36.942 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 55.873 36.987 55.907 ;
      VIA 36.942 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 55.333 36.987 55.367 ;
      VIA 36.942 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 54.793 36.987 54.827 ;
      VIA 36.942 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 54.253 36.987 54.287 ;
      VIA 36.942 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 53.713 36.987 53.747 ;
      VIA 36.942 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 53.173 36.987 53.207 ;
      VIA 36.942 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 52.633 36.987 52.667 ;
      VIA 36.942 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 52.093 36.987 52.127 ;
      VIA 36.942 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 51.553 36.987 51.587 ;
      VIA 36.942 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 51.013 36.987 51.047 ;
      VIA 36.942 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 50.473 36.987 50.507 ;
      VIA 36.942 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 49.933 36.987 49.967 ;
      VIA 36.942 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 49.393 36.987 49.427 ;
      VIA 36.942 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 48.853 36.987 48.887 ;
      VIA 36.942 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 48.313 36.987 48.347 ;
      VIA 36.942 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 47.773 36.987 47.807 ;
      VIA 36.942 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 47.233 36.987 47.267 ;
      VIA 36.942 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 46.693 36.987 46.727 ;
      VIA 36.942 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 46.153 36.987 46.187 ;
      VIA 36.942 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 45.613 36.987 45.647 ;
      VIA 36.942 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 45.073 36.987 45.107 ;
      VIA 36.942 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 44.533 36.987 44.567 ;
      VIA 36.942 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 43.993 36.987 44.027 ;
      VIA 36.942 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 43.453 36.987 43.487 ;
      VIA 36.942 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 42.913 36.987 42.947 ;
      VIA 36.942 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 42.373 36.987 42.407 ;
      VIA 36.942 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 41.833 36.987 41.867 ;
      VIA 36.942 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 41.293 36.987 41.327 ;
      VIA 36.942 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 40.753 36.987 40.787 ;
      VIA 36.942 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 40.213 36.987 40.247 ;
      VIA 36.942 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.673 36.987 39.707 ;
      VIA 36.942 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.133 36.987 39.167 ;
      VIA 36.942 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.593 36.987 38.627 ;
      VIA 36.942 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.053 36.987 38.087 ;
      VIA 36.942 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 37.513 36.987 37.547 ;
      VIA 36.942 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.973 36.987 37.007 ;
      VIA 36.942 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.433 36.987 36.467 ;
      VIA 36.942 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.893 36.987 35.927 ;
      VIA 36.942 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.353 36.987 35.387 ;
      VIA 36.942 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.813 36.987 34.847 ;
      VIA 36.942 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.273 36.987 34.307 ;
      VIA 36.942 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.733 36.987 33.767 ;
      VIA 36.942 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.193 36.987 33.227 ;
      VIA 36.942 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.653 36.987 32.687 ;
      VIA 36.942 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.113 36.987 32.147 ;
      VIA 36.942 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.573 36.987 31.607 ;
      VIA 36.942 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.033 36.987 31.067 ;
      VIA 36.942 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 30.493 36.987 30.527 ;
      VIA 36.942 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.953 36.987 29.987 ;
      VIA 36.942 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.413 36.987 29.447 ;
      VIA 36.942 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.873 36.987 28.907 ;
      VIA 36.942 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.333 36.987 28.367 ;
      VIA 36.942 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.793 36.987 27.827 ;
      VIA 36.942 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.253 36.987 27.287 ;
      VIA 36.942 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.713 36.987 26.747 ;
      VIA 36.942 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.173 36.987 26.207 ;
      VIA 36.942 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.633 36.987 25.667 ;
      VIA 36.942 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.093 36.987 25.127 ;
      VIA 36.942 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.553 36.987 24.587 ;
      VIA 36.942 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.013 36.987 24.047 ;
      VIA 36.942 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 23.473 36.987 23.507 ;
      VIA 36.942 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.933 36.987 22.967 ;
      VIA 36.942 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.393 36.987 22.427 ;
      VIA 36.942 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.853 36.987 21.887 ;
      VIA 36.942 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.313 36.987 21.347 ;
      VIA 36.942 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.773 36.987 20.807 ;
      VIA 36.942 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.233 36.987 20.267 ;
      VIA 36.942 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.693 36.987 19.727 ;
      VIA 36.942 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.153 36.987 19.187 ;
      VIA 36.942 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.613 36.987 18.647 ;
      VIA 36.942 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.073 36.987 18.107 ;
      VIA 36.942 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 17.533 36.987 17.567 ;
      VIA 36.942 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.993 36.987 17.027 ;
      VIA 36.942 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.453 36.987 16.487 ;
      VIA 36.942 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.913 36.987 15.947 ;
      VIA 36.942 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.373 36.987 15.407 ;
      VIA 36.942 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.833 36.987 14.867 ;
      VIA 36.942 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.293 36.987 14.327 ;
      VIA 36.942 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.753 36.987 13.787 ;
      VIA 36.942 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.213 36.987 13.247 ;
      VIA 36.942 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.673 36.987 12.707 ;
      VIA 36.942 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.133 36.987 12.167 ;
      VIA 36.942 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.593 36.987 11.627 ;
      VIA 36.942 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.053 36.987 11.087 ;
      VIA 36.942 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 10.513 36.987 10.547 ;
      VIA 36.942 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.973 36.987 10.007 ;
      VIA 36.942 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.433 36.987 9.467 ;
      VIA 36.942 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.893 36.987 8.927 ;
      VIA 36.942 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.353 36.987 8.387 ;
      VIA 36.942 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.813 36.987 7.847 ;
      VIA 36.942 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.273 36.987 7.307 ;
      VIA 36.942 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.733 36.987 6.767 ;
      VIA 36.942 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.193 36.987 6.227 ;
      VIA 36.942 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.653 36.987 5.687 ;
      VIA 36.942 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.113 36.987 5.147 ;
      VIA 36.942 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.573 36.987 4.607 ;
      VIA 36.942 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.033 36.987 4.067 ;
      VIA 36.942 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 3.493 36.987 3.527 ;
      VIA 36.942 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.953 36.987 2.987 ;
      VIA 36.942 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.413 36.987 2.447 ;
      VIA 36.942 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.873 36.987 1.907 ;
      VIA 36.942 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.333 36.987 1.367 ;
      VIA 36.942 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 73.153 31.083 73.187 ;
      VIA 31.038 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 72.613 31.083 72.647 ;
      VIA 31.038 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 72.073 31.083 72.107 ;
      VIA 31.038 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 71.533 31.083 71.567 ;
      VIA 31.038 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 70.993 31.083 71.027 ;
      VIA 31.038 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 70.453 31.083 70.487 ;
      VIA 31.038 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 69.913 31.083 69.947 ;
      VIA 31.038 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 69.373 31.083 69.407 ;
      VIA 31.038 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 68.833 31.083 68.867 ;
      VIA 31.038 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 68.293 31.083 68.327 ;
      VIA 31.038 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 67.753 31.083 67.787 ;
      VIA 31.038 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 67.213 31.083 67.247 ;
      VIA 31.038 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 66.673 31.083 66.707 ;
      VIA 31.038 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 66.133 31.083 66.167 ;
      VIA 31.038 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 65.593 31.083 65.627 ;
      VIA 31.038 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 65.053 31.083 65.087 ;
      VIA 31.038 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 64.513 31.083 64.547 ;
      VIA 31.038 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 63.973 31.083 64.007 ;
      VIA 31.038 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 63.433 31.083 63.467 ;
      VIA 31.038 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 62.893 31.083 62.927 ;
      VIA 31.038 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 62.353 31.083 62.387 ;
      VIA 31.038 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 61.813 31.083 61.847 ;
      VIA 31.038 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 61.273 31.083 61.307 ;
      VIA 31.038 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 60.733 31.083 60.767 ;
      VIA 31.038 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 60.193 31.083 60.227 ;
      VIA 31.038 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 59.653 31.083 59.687 ;
      VIA 31.038 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 59.113 31.083 59.147 ;
      VIA 31.038 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 58.573 31.083 58.607 ;
      VIA 31.038 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 58.033 31.083 58.067 ;
      VIA 31.038 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 57.493 31.083 57.527 ;
      VIA 31.038 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 56.953 31.083 56.987 ;
      VIA 31.038 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 56.413 31.083 56.447 ;
      VIA 31.038 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 55.873 31.083 55.907 ;
      VIA 31.038 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 55.333 31.083 55.367 ;
      VIA 31.038 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 54.793 31.083 54.827 ;
      VIA 31.038 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 54.253 31.083 54.287 ;
      VIA 31.038 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 53.713 31.083 53.747 ;
      VIA 31.038 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 53.173 31.083 53.207 ;
      VIA 31.038 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 52.633 31.083 52.667 ;
      VIA 31.038 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 52.093 31.083 52.127 ;
      VIA 31.038 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 51.553 31.083 51.587 ;
      VIA 31.038 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 51.013 31.083 51.047 ;
      VIA 31.038 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 50.473 31.083 50.507 ;
      VIA 31.038 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 49.933 31.083 49.967 ;
      VIA 31.038 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 49.393 31.083 49.427 ;
      VIA 31.038 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 48.853 31.083 48.887 ;
      VIA 31.038 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 48.313 31.083 48.347 ;
      VIA 31.038 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 47.773 31.083 47.807 ;
      VIA 31.038 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 47.233 31.083 47.267 ;
      VIA 31.038 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 46.693 31.083 46.727 ;
      VIA 31.038 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 46.153 31.083 46.187 ;
      VIA 31.038 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 45.613 31.083 45.647 ;
      VIA 31.038 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 45.073 31.083 45.107 ;
      VIA 31.038 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 44.533 31.083 44.567 ;
      VIA 31.038 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 43.993 31.083 44.027 ;
      VIA 31.038 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 43.453 31.083 43.487 ;
      VIA 31.038 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 42.913 31.083 42.947 ;
      VIA 31.038 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 42.373 31.083 42.407 ;
      VIA 31.038 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 41.833 31.083 41.867 ;
      VIA 31.038 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 41.293 31.083 41.327 ;
      VIA 31.038 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 40.753 31.083 40.787 ;
      VIA 31.038 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 40.213 31.083 40.247 ;
      VIA 31.038 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.673 31.083 39.707 ;
      VIA 31.038 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.133 31.083 39.167 ;
      VIA 31.038 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.593 31.083 38.627 ;
      VIA 31.038 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.053 31.083 38.087 ;
      VIA 31.038 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 37.513 31.083 37.547 ;
      VIA 31.038 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.973 31.083 37.007 ;
      VIA 31.038 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.433 31.083 36.467 ;
      VIA 31.038 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.893 31.083 35.927 ;
      VIA 31.038 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.353 31.083 35.387 ;
      VIA 31.038 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.813 31.083 34.847 ;
      VIA 31.038 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.273 31.083 34.307 ;
      VIA 31.038 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.733 31.083 33.767 ;
      VIA 31.038 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.193 31.083 33.227 ;
      VIA 31.038 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.653 31.083 32.687 ;
      VIA 31.038 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.113 31.083 32.147 ;
      VIA 31.038 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.573 31.083 31.607 ;
      VIA 31.038 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.033 31.083 31.067 ;
      VIA 31.038 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 30.493 31.083 30.527 ;
      VIA 31.038 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.953 31.083 29.987 ;
      VIA 31.038 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.413 31.083 29.447 ;
      VIA 31.038 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.873 31.083 28.907 ;
      VIA 31.038 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.333 31.083 28.367 ;
      VIA 31.038 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.793 31.083 27.827 ;
      VIA 31.038 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.253 31.083 27.287 ;
      VIA 31.038 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.713 31.083 26.747 ;
      VIA 31.038 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.173 31.083 26.207 ;
      VIA 31.038 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.633 31.083 25.667 ;
      VIA 31.038 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.093 31.083 25.127 ;
      VIA 31.038 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.553 31.083 24.587 ;
      VIA 31.038 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.013 31.083 24.047 ;
      VIA 31.038 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 23.473 31.083 23.507 ;
      VIA 31.038 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.933 31.083 22.967 ;
      VIA 31.038 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.393 31.083 22.427 ;
      VIA 31.038 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.853 31.083 21.887 ;
      VIA 31.038 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.313 31.083 21.347 ;
      VIA 31.038 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.773 31.083 20.807 ;
      VIA 31.038 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.233 31.083 20.267 ;
      VIA 31.038 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.693 31.083 19.727 ;
      VIA 31.038 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.153 31.083 19.187 ;
      VIA 31.038 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.613 31.083 18.647 ;
      VIA 31.038 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.073 31.083 18.107 ;
      VIA 31.038 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 17.533 31.083 17.567 ;
      VIA 31.038 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.993 31.083 17.027 ;
      VIA 31.038 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.453 31.083 16.487 ;
      VIA 31.038 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.913 31.083 15.947 ;
      VIA 31.038 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.373 31.083 15.407 ;
      VIA 31.038 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.833 31.083 14.867 ;
      VIA 31.038 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.293 31.083 14.327 ;
      VIA 31.038 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.753 31.083 13.787 ;
      VIA 31.038 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.213 31.083 13.247 ;
      VIA 31.038 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.673 31.083 12.707 ;
      VIA 31.038 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.133 31.083 12.167 ;
      VIA 31.038 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.593 31.083 11.627 ;
      VIA 31.038 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.053 31.083 11.087 ;
      VIA 31.038 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 10.513 31.083 10.547 ;
      VIA 31.038 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.973 31.083 10.007 ;
      VIA 31.038 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.433 31.083 9.467 ;
      VIA 31.038 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.893 31.083 8.927 ;
      VIA 31.038 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.353 31.083 8.387 ;
      VIA 31.038 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.813 31.083 7.847 ;
      VIA 31.038 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.273 31.083 7.307 ;
      VIA 31.038 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.733 31.083 6.767 ;
      VIA 31.038 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.193 31.083 6.227 ;
      VIA 31.038 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.653 31.083 5.687 ;
      VIA 31.038 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.113 31.083 5.147 ;
      VIA 31.038 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.573 31.083 4.607 ;
      VIA 31.038 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.033 31.083 4.067 ;
      VIA 31.038 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 3.493 31.083 3.527 ;
      VIA 31.038 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.953 31.083 2.987 ;
      VIA 31.038 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.413 31.083 2.447 ;
      VIA 31.038 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.873 31.083 1.907 ;
      VIA 31.038 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.333 31.083 1.367 ;
      VIA 31.038 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 73.153 25.179 73.187 ;
      VIA 25.134 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 72.613 25.179 72.647 ;
      VIA 25.134 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 72.073 25.179 72.107 ;
      VIA 25.134 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 71.533 25.179 71.567 ;
      VIA 25.134 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 70.993 25.179 71.027 ;
      VIA 25.134 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 70.453 25.179 70.487 ;
      VIA 25.134 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 69.913 25.179 69.947 ;
      VIA 25.134 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 69.373 25.179 69.407 ;
      VIA 25.134 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 68.833 25.179 68.867 ;
      VIA 25.134 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 68.293 25.179 68.327 ;
      VIA 25.134 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 67.753 25.179 67.787 ;
      VIA 25.134 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 67.213 25.179 67.247 ;
      VIA 25.134 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 66.673 25.179 66.707 ;
      VIA 25.134 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 66.133 25.179 66.167 ;
      VIA 25.134 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 65.593 25.179 65.627 ;
      VIA 25.134 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 65.053 25.179 65.087 ;
      VIA 25.134 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 64.513 25.179 64.547 ;
      VIA 25.134 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 63.973 25.179 64.007 ;
      VIA 25.134 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 63.433 25.179 63.467 ;
      VIA 25.134 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 62.893 25.179 62.927 ;
      VIA 25.134 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 62.353 25.179 62.387 ;
      VIA 25.134 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 61.813 25.179 61.847 ;
      VIA 25.134 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 61.273 25.179 61.307 ;
      VIA 25.134 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 60.733 25.179 60.767 ;
      VIA 25.134 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 60.193 25.179 60.227 ;
      VIA 25.134 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 59.653 25.179 59.687 ;
      VIA 25.134 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 59.113 25.179 59.147 ;
      VIA 25.134 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 58.573 25.179 58.607 ;
      VIA 25.134 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 58.033 25.179 58.067 ;
      VIA 25.134 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 57.493 25.179 57.527 ;
      VIA 25.134 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 56.953 25.179 56.987 ;
      VIA 25.134 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 56.413 25.179 56.447 ;
      VIA 25.134 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 55.873 25.179 55.907 ;
      VIA 25.134 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 55.333 25.179 55.367 ;
      VIA 25.134 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 54.793 25.179 54.827 ;
      VIA 25.134 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 54.253 25.179 54.287 ;
      VIA 25.134 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 53.713 25.179 53.747 ;
      VIA 25.134 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 53.173 25.179 53.207 ;
      VIA 25.134 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 52.633 25.179 52.667 ;
      VIA 25.134 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 52.093 25.179 52.127 ;
      VIA 25.134 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 51.553 25.179 51.587 ;
      VIA 25.134 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 51.013 25.179 51.047 ;
      VIA 25.134 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 50.473 25.179 50.507 ;
      VIA 25.134 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 49.933 25.179 49.967 ;
      VIA 25.134 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 49.393 25.179 49.427 ;
      VIA 25.134 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 48.853 25.179 48.887 ;
      VIA 25.134 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 48.313 25.179 48.347 ;
      VIA 25.134 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 47.773 25.179 47.807 ;
      VIA 25.134 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 47.233 25.179 47.267 ;
      VIA 25.134 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 46.693 25.179 46.727 ;
      VIA 25.134 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 46.153 25.179 46.187 ;
      VIA 25.134 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 45.613 25.179 45.647 ;
      VIA 25.134 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 45.073 25.179 45.107 ;
      VIA 25.134 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 44.533 25.179 44.567 ;
      VIA 25.134 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 43.993 25.179 44.027 ;
      VIA 25.134 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 43.453 25.179 43.487 ;
      VIA 25.134 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 42.913 25.179 42.947 ;
      VIA 25.134 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 42.373 25.179 42.407 ;
      VIA 25.134 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 41.833 25.179 41.867 ;
      VIA 25.134 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 41.293 25.179 41.327 ;
      VIA 25.134 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 40.753 25.179 40.787 ;
      VIA 25.134 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 40.213 25.179 40.247 ;
      VIA 25.134 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.673 25.179 39.707 ;
      VIA 25.134 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.133 25.179 39.167 ;
      VIA 25.134 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.593 25.179 38.627 ;
      VIA 25.134 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.053 25.179 38.087 ;
      VIA 25.134 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 37.513 25.179 37.547 ;
      VIA 25.134 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.973 25.179 37.007 ;
      VIA 25.134 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.433 25.179 36.467 ;
      VIA 25.134 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.893 25.179 35.927 ;
      VIA 25.134 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.353 25.179 35.387 ;
      VIA 25.134 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.813 25.179 34.847 ;
      VIA 25.134 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.273 25.179 34.307 ;
      VIA 25.134 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.733 25.179 33.767 ;
      VIA 25.134 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.193 25.179 33.227 ;
      VIA 25.134 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.653 25.179 32.687 ;
      VIA 25.134 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.113 25.179 32.147 ;
      VIA 25.134 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.573 25.179 31.607 ;
      VIA 25.134 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.033 25.179 31.067 ;
      VIA 25.134 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 30.493 25.179 30.527 ;
      VIA 25.134 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.953 25.179 29.987 ;
      VIA 25.134 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.413 25.179 29.447 ;
      VIA 25.134 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.873 25.179 28.907 ;
      VIA 25.134 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.333 25.179 28.367 ;
      VIA 25.134 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.793 25.179 27.827 ;
      VIA 25.134 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.253 25.179 27.287 ;
      VIA 25.134 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.713 25.179 26.747 ;
      VIA 25.134 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.173 25.179 26.207 ;
      VIA 25.134 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.633 25.179 25.667 ;
      VIA 25.134 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.093 25.179 25.127 ;
      VIA 25.134 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.553 25.179 24.587 ;
      VIA 25.134 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.013 25.179 24.047 ;
      VIA 25.134 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 23.473 25.179 23.507 ;
      VIA 25.134 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.933 25.179 22.967 ;
      VIA 25.134 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.393 25.179 22.427 ;
      VIA 25.134 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.853 25.179 21.887 ;
      VIA 25.134 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.313 25.179 21.347 ;
      VIA 25.134 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.773 25.179 20.807 ;
      VIA 25.134 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.233 25.179 20.267 ;
      VIA 25.134 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.693 25.179 19.727 ;
      VIA 25.134 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.153 25.179 19.187 ;
      VIA 25.134 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.613 25.179 18.647 ;
      VIA 25.134 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.073 25.179 18.107 ;
      VIA 25.134 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 17.533 25.179 17.567 ;
      VIA 25.134 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.993 25.179 17.027 ;
      VIA 25.134 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.453 25.179 16.487 ;
      VIA 25.134 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.913 25.179 15.947 ;
      VIA 25.134 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.373 25.179 15.407 ;
      VIA 25.134 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.833 25.179 14.867 ;
      VIA 25.134 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.293 25.179 14.327 ;
      VIA 25.134 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.753 25.179 13.787 ;
      VIA 25.134 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.213 25.179 13.247 ;
      VIA 25.134 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.673 25.179 12.707 ;
      VIA 25.134 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.133 25.179 12.167 ;
      VIA 25.134 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.593 25.179 11.627 ;
      VIA 25.134 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.053 25.179 11.087 ;
      VIA 25.134 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 10.513 25.179 10.547 ;
      VIA 25.134 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.973 25.179 10.007 ;
      VIA 25.134 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.433 25.179 9.467 ;
      VIA 25.134 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.893 25.179 8.927 ;
      VIA 25.134 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.353 25.179 8.387 ;
      VIA 25.134 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.813 25.179 7.847 ;
      VIA 25.134 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.273 25.179 7.307 ;
      VIA 25.134 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.733 25.179 6.767 ;
      VIA 25.134 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.193 25.179 6.227 ;
      VIA 25.134 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.653 25.179 5.687 ;
      VIA 25.134 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.113 25.179 5.147 ;
      VIA 25.134 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.573 25.179 4.607 ;
      VIA 25.134 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.033 25.179 4.067 ;
      VIA 25.134 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 3.493 25.179 3.527 ;
      VIA 25.134 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.953 25.179 2.987 ;
      VIA 25.134 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.413 25.179 2.447 ;
      VIA 25.134 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.873 25.179 1.907 ;
      VIA 25.134 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.333 25.179 1.367 ;
      VIA 25.134 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 73.153 19.275 73.187 ;
      VIA 19.23 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 72.613 19.275 72.647 ;
      VIA 19.23 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 72.073 19.275 72.107 ;
      VIA 19.23 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 71.533 19.275 71.567 ;
      VIA 19.23 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 70.993 19.275 71.027 ;
      VIA 19.23 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 70.453 19.275 70.487 ;
      VIA 19.23 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 69.913 19.275 69.947 ;
      VIA 19.23 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 69.373 19.275 69.407 ;
      VIA 19.23 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 68.833 19.275 68.867 ;
      VIA 19.23 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 68.293 19.275 68.327 ;
      VIA 19.23 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 67.753 19.275 67.787 ;
      VIA 19.23 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 67.213 19.275 67.247 ;
      VIA 19.23 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 66.673 19.275 66.707 ;
      VIA 19.23 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 66.133 19.275 66.167 ;
      VIA 19.23 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 65.593 19.275 65.627 ;
      VIA 19.23 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 65.053 19.275 65.087 ;
      VIA 19.23 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 64.513 19.275 64.547 ;
      VIA 19.23 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 63.973 19.275 64.007 ;
      VIA 19.23 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 63.433 19.275 63.467 ;
      VIA 19.23 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 62.893 19.275 62.927 ;
      VIA 19.23 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 62.353 19.275 62.387 ;
      VIA 19.23 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 61.813 19.275 61.847 ;
      VIA 19.23 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 61.273 19.275 61.307 ;
      VIA 19.23 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 60.733 19.275 60.767 ;
      VIA 19.23 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 60.193 19.275 60.227 ;
      VIA 19.23 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 59.653 19.275 59.687 ;
      VIA 19.23 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 59.113 19.275 59.147 ;
      VIA 19.23 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 58.573 19.275 58.607 ;
      VIA 19.23 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 58.033 19.275 58.067 ;
      VIA 19.23 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 57.493 19.275 57.527 ;
      VIA 19.23 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 56.953 19.275 56.987 ;
      VIA 19.23 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 56.413 19.275 56.447 ;
      VIA 19.23 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 55.873 19.275 55.907 ;
      VIA 19.23 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 55.333 19.275 55.367 ;
      VIA 19.23 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 54.793 19.275 54.827 ;
      VIA 19.23 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 54.253 19.275 54.287 ;
      VIA 19.23 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 53.713 19.275 53.747 ;
      VIA 19.23 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 53.173 19.275 53.207 ;
      VIA 19.23 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 52.633 19.275 52.667 ;
      VIA 19.23 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 52.093 19.275 52.127 ;
      VIA 19.23 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 51.553 19.275 51.587 ;
      VIA 19.23 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 51.013 19.275 51.047 ;
      VIA 19.23 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 50.473 19.275 50.507 ;
      VIA 19.23 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 49.933 19.275 49.967 ;
      VIA 19.23 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 49.393 19.275 49.427 ;
      VIA 19.23 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 48.853 19.275 48.887 ;
      VIA 19.23 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 48.313 19.275 48.347 ;
      VIA 19.23 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 47.773 19.275 47.807 ;
      VIA 19.23 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 47.233 19.275 47.267 ;
      VIA 19.23 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 46.693 19.275 46.727 ;
      VIA 19.23 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 46.153 19.275 46.187 ;
      VIA 19.23 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 45.613 19.275 45.647 ;
      VIA 19.23 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 45.073 19.275 45.107 ;
      VIA 19.23 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 44.533 19.275 44.567 ;
      VIA 19.23 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 43.993 19.275 44.027 ;
      VIA 19.23 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 43.453 19.275 43.487 ;
      VIA 19.23 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 42.913 19.275 42.947 ;
      VIA 19.23 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 42.373 19.275 42.407 ;
      VIA 19.23 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 41.833 19.275 41.867 ;
      VIA 19.23 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 41.293 19.275 41.327 ;
      VIA 19.23 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 40.753 19.275 40.787 ;
      VIA 19.23 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 40.213 19.275 40.247 ;
      VIA 19.23 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.673 19.275 39.707 ;
      VIA 19.23 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.133 19.275 39.167 ;
      VIA 19.23 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.593 19.275 38.627 ;
      VIA 19.23 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.053 19.275 38.087 ;
      VIA 19.23 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 37.513 19.275 37.547 ;
      VIA 19.23 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.973 19.275 37.007 ;
      VIA 19.23 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.433 19.275 36.467 ;
      VIA 19.23 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.893 19.275 35.927 ;
      VIA 19.23 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.353 19.275 35.387 ;
      VIA 19.23 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.813 19.275 34.847 ;
      VIA 19.23 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.273 19.275 34.307 ;
      VIA 19.23 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.733 19.275 33.767 ;
      VIA 19.23 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.193 19.275 33.227 ;
      VIA 19.23 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.653 19.275 32.687 ;
      VIA 19.23 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.113 19.275 32.147 ;
      VIA 19.23 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.573 19.275 31.607 ;
      VIA 19.23 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.033 19.275 31.067 ;
      VIA 19.23 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 30.493 19.275 30.527 ;
      VIA 19.23 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.953 19.275 29.987 ;
      VIA 19.23 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.413 19.275 29.447 ;
      VIA 19.23 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.873 19.275 28.907 ;
      VIA 19.23 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.333 19.275 28.367 ;
      VIA 19.23 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.793 19.275 27.827 ;
      VIA 19.23 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.253 19.275 27.287 ;
      VIA 19.23 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.713 19.275 26.747 ;
      VIA 19.23 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.173 19.275 26.207 ;
      VIA 19.23 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.633 19.275 25.667 ;
      VIA 19.23 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.093 19.275 25.127 ;
      VIA 19.23 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.553 19.275 24.587 ;
      VIA 19.23 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.013 19.275 24.047 ;
      VIA 19.23 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 23.473 19.275 23.507 ;
      VIA 19.23 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.933 19.275 22.967 ;
      VIA 19.23 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.393 19.275 22.427 ;
      VIA 19.23 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.853 19.275 21.887 ;
      VIA 19.23 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.313 19.275 21.347 ;
      VIA 19.23 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.773 19.275 20.807 ;
      VIA 19.23 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.233 19.275 20.267 ;
      VIA 19.23 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.693 19.275 19.727 ;
      VIA 19.23 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.153 19.275 19.187 ;
      VIA 19.23 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.613 19.275 18.647 ;
      VIA 19.23 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.073 19.275 18.107 ;
      VIA 19.23 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 17.533 19.275 17.567 ;
      VIA 19.23 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.993 19.275 17.027 ;
      VIA 19.23 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.453 19.275 16.487 ;
      VIA 19.23 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.913 19.275 15.947 ;
      VIA 19.23 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.373 19.275 15.407 ;
      VIA 19.23 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.833 19.275 14.867 ;
      VIA 19.23 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.293 19.275 14.327 ;
      VIA 19.23 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.753 19.275 13.787 ;
      VIA 19.23 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.213 19.275 13.247 ;
      VIA 19.23 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.673 19.275 12.707 ;
      VIA 19.23 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.133 19.275 12.167 ;
      VIA 19.23 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.593 19.275 11.627 ;
      VIA 19.23 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.053 19.275 11.087 ;
      VIA 19.23 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 10.513 19.275 10.547 ;
      VIA 19.23 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.973 19.275 10.007 ;
      VIA 19.23 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.433 19.275 9.467 ;
      VIA 19.23 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.893 19.275 8.927 ;
      VIA 19.23 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.353 19.275 8.387 ;
      VIA 19.23 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.813 19.275 7.847 ;
      VIA 19.23 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.273 19.275 7.307 ;
      VIA 19.23 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.733 19.275 6.767 ;
      VIA 19.23 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.193 19.275 6.227 ;
      VIA 19.23 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.653 19.275 5.687 ;
      VIA 19.23 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.113 19.275 5.147 ;
      VIA 19.23 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.573 19.275 4.607 ;
      VIA 19.23 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.033 19.275 4.067 ;
      VIA 19.23 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 3.493 19.275 3.527 ;
      VIA 19.23 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.953 19.275 2.987 ;
      VIA 19.23 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.413 19.275 2.447 ;
      VIA 19.23 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.873 19.275 1.907 ;
      VIA 19.23 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.333 19.275 1.367 ;
      VIA 19.23 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 73.153 13.371 73.187 ;
      VIA 13.326 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 72.613 13.371 72.647 ;
      VIA 13.326 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 72.073 13.371 72.107 ;
      VIA 13.326 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 71.533 13.371 71.567 ;
      VIA 13.326 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 70.993 13.371 71.027 ;
      VIA 13.326 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 70.453 13.371 70.487 ;
      VIA 13.326 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 69.913 13.371 69.947 ;
      VIA 13.326 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 69.373 13.371 69.407 ;
      VIA 13.326 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 68.833 13.371 68.867 ;
      VIA 13.326 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 68.293 13.371 68.327 ;
      VIA 13.326 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 67.753 13.371 67.787 ;
      VIA 13.326 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 67.213 13.371 67.247 ;
      VIA 13.326 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 66.673 13.371 66.707 ;
      VIA 13.326 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 66.133 13.371 66.167 ;
      VIA 13.326 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 65.593 13.371 65.627 ;
      VIA 13.326 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 65.053 13.371 65.087 ;
      VIA 13.326 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 64.513 13.371 64.547 ;
      VIA 13.326 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 63.973 13.371 64.007 ;
      VIA 13.326 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 63.433 13.371 63.467 ;
      VIA 13.326 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 62.893 13.371 62.927 ;
      VIA 13.326 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 62.353 13.371 62.387 ;
      VIA 13.326 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 61.813 13.371 61.847 ;
      VIA 13.326 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 61.273 13.371 61.307 ;
      VIA 13.326 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 60.733 13.371 60.767 ;
      VIA 13.326 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 60.193 13.371 60.227 ;
      VIA 13.326 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 59.653 13.371 59.687 ;
      VIA 13.326 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 59.113 13.371 59.147 ;
      VIA 13.326 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 58.573 13.371 58.607 ;
      VIA 13.326 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 58.033 13.371 58.067 ;
      VIA 13.326 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 57.493 13.371 57.527 ;
      VIA 13.326 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 56.953 13.371 56.987 ;
      VIA 13.326 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 56.413 13.371 56.447 ;
      VIA 13.326 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 55.873 13.371 55.907 ;
      VIA 13.326 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 55.333 13.371 55.367 ;
      VIA 13.326 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 54.793 13.371 54.827 ;
      VIA 13.326 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 54.253 13.371 54.287 ;
      VIA 13.326 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 53.713 13.371 53.747 ;
      VIA 13.326 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 53.173 13.371 53.207 ;
      VIA 13.326 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 52.633 13.371 52.667 ;
      VIA 13.326 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 52.093 13.371 52.127 ;
      VIA 13.326 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 51.553 13.371 51.587 ;
      VIA 13.326 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 51.013 13.371 51.047 ;
      VIA 13.326 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 50.473 13.371 50.507 ;
      VIA 13.326 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 49.933 13.371 49.967 ;
      VIA 13.326 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 49.393 13.371 49.427 ;
      VIA 13.326 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 48.853 13.371 48.887 ;
      VIA 13.326 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 48.313 13.371 48.347 ;
      VIA 13.326 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 47.773 13.371 47.807 ;
      VIA 13.326 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 47.233 13.371 47.267 ;
      VIA 13.326 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 46.693 13.371 46.727 ;
      VIA 13.326 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 46.153 13.371 46.187 ;
      VIA 13.326 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 45.613 13.371 45.647 ;
      VIA 13.326 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 45.073 13.371 45.107 ;
      VIA 13.326 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 44.533 13.371 44.567 ;
      VIA 13.326 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 43.993 13.371 44.027 ;
      VIA 13.326 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 43.453 13.371 43.487 ;
      VIA 13.326 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 42.913 13.371 42.947 ;
      VIA 13.326 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 42.373 13.371 42.407 ;
      VIA 13.326 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 41.833 13.371 41.867 ;
      VIA 13.326 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 41.293 13.371 41.327 ;
      VIA 13.326 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 40.753 13.371 40.787 ;
      VIA 13.326 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 40.213 13.371 40.247 ;
      VIA 13.326 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.673 13.371 39.707 ;
      VIA 13.326 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.133 13.371 39.167 ;
      VIA 13.326 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.593 13.371 38.627 ;
      VIA 13.326 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.053 13.371 38.087 ;
      VIA 13.326 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 37.513 13.371 37.547 ;
      VIA 13.326 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.973 13.371 37.007 ;
      VIA 13.326 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.433 13.371 36.467 ;
      VIA 13.326 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.893 13.371 35.927 ;
      VIA 13.326 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.353 13.371 35.387 ;
      VIA 13.326 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.813 13.371 34.847 ;
      VIA 13.326 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.273 13.371 34.307 ;
      VIA 13.326 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.733 13.371 33.767 ;
      VIA 13.326 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.193 13.371 33.227 ;
      VIA 13.326 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.653 13.371 32.687 ;
      VIA 13.326 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.113 13.371 32.147 ;
      VIA 13.326 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.573 13.371 31.607 ;
      VIA 13.326 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.033 13.371 31.067 ;
      VIA 13.326 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 30.493 13.371 30.527 ;
      VIA 13.326 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.953 13.371 29.987 ;
      VIA 13.326 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.413 13.371 29.447 ;
      VIA 13.326 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.873 13.371 28.907 ;
      VIA 13.326 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.333 13.371 28.367 ;
      VIA 13.326 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.793 13.371 27.827 ;
      VIA 13.326 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.253 13.371 27.287 ;
      VIA 13.326 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.713 13.371 26.747 ;
      VIA 13.326 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.173 13.371 26.207 ;
      VIA 13.326 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.633 13.371 25.667 ;
      VIA 13.326 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.093 13.371 25.127 ;
      VIA 13.326 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.553 13.371 24.587 ;
      VIA 13.326 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.013 13.371 24.047 ;
      VIA 13.326 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 23.473 13.371 23.507 ;
      VIA 13.326 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.933 13.371 22.967 ;
      VIA 13.326 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.393 13.371 22.427 ;
      VIA 13.326 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.853 13.371 21.887 ;
      VIA 13.326 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.313 13.371 21.347 ;
      VIA 13.326 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.773 13.371 20.807 ;
      VIA 13.326 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.233 13.371 20.267 ;
      VIA 13.326 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.693 13.371 19.727 ;
      VIA 13.326 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.153 13.371 19.187 ;
      VIA 13.326 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.613 13.371 18.647 ;
      VIA 13.326 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.073 13.371 18.107 ;
      VIA 13.326 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 17.533 13.371 17.567 ;
      VIA 13.326 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.993 13.371 17.027 ;
      VIA 13.326 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.453 13.371 16.487 ;
      VIA 13.326 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.913 13.371 15.947 ;
      VIA 13.326 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.373 13.371 15.407 ;
      VIA 13.326 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.833 13.371 14.867 ;
      VIA 13.326 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.293 13.371 14.327 ;
      VIA 13.326 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.753 13.371 13.787 ;
      VIA 13.326 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.213 13.371 13.247 ;
      VIA 13.326 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.673 13.371 12.707 ;
      VIA 13.326 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.133 13.371 12.167 ;
      VIA 13.326 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.593 13.371 11.627 ;
      VIA 13.326 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.053 13.371 11.087 ;
      VIA 13.326 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 10.513 13.371 10.547 ;
      VIA 13.326 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.973 13.371 10.007 ;
      VIA 13.326 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.433 13.371 9.467 ;
      VIA 13.326 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.893 13.371 8.927 ;
      VIA 13.326 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.353 13.371 8.387 ;
      VIA 13.326 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.813 13.371 7.847 ;
      VIA 13.326 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.273 13.371 7.307 ;
      VIA 13.326 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.733 13.371 6.767 ;
      VIA 13.326 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.193 13.371 6.227 ;
      VIA 13.326 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.653 13.371 5.687 ;
      VIA 13.326 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.113 13.371 5.147 ;
      VIA 13.326 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.573 13.371 4.607 ;
      VIA 13.326 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.033 13.371 4.067 ;
      VIA 13.326 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 3.493 13.371 3.527 ;
      VIA 13.326 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.953 13.371 2.987 ;
      VIA 13.326 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.413 13.371 2.447 ;
      VIA 13.326 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.873 13.371 1.907 ;
      VIA 13.326 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.333 13.371 1.367 ;
      VIA 13.326 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 73.153 7.467 73.187 ;
      VIA 7.422 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 72.613 7.467 72.647 ;
      VIA 7.422 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 72.073 7.467 72.107 ;
      VIA 7.422 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 71.533 7.467 71.567 ;
      VIA 7.422 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 70.993 7.467 71.027 ;
      VIA 7.422 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 70.453 7.467 70.487 ;
      VIA 7.422 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 69.913 7.467 69.947 ;
      VIA 7.422 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 69.373 7.467 69.407 ;
      VIA 7.422 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 68.833 7.467 68.867 ;
      VIA 7.422 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 68.293 7.467 68.327 ;
      VIA 7.422 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 67.753 7.467 67.787 ;
      VIA 7.422 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 67.213 7.467 67.247 ;
      VIA 7.422 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 66.673 7.467 66.707 ;
      VIA 7.422 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 66.133 7.467 66.167 ;
      VIA 7.422 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 65.593 7.467 65.627 ;
      VIA 7.422 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 65.053 7.467 65.087 ;
      VIA 7.422 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 64.513 7.467 64.547 ;
      VIA 7.422 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 63.973 7.467 64.007 ;
      VIA 7.422 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 63.433 7.467 63.467 ;
      VIA 7.422 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 62.893 7.467 62.927 ;
      VIA 7.422 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 62.353 7.467 62.387 ;
      VIA 7.422 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 61.813 7.467 61.847 ;
      VIA 7.422 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 61.273 7.467 61.307 ;
      VIA 7.422 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 60.733 7.467 60.767 ;
      VIA 7.422 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 60.193 7.467 60.227 ;
      VIA 7.422 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 59.653 7.467 59.687 ;
      VIA 7.422 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 59.113 7.467 59.147 ;
      VIA 7.422 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 58.573 7.467 58.607 ;
      VIA 7.422 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 58.033 7.467 58.067 ;
      VIA 7.422 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 57.493 7.467 57.527 ;
      VIA 7.422 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 56.953 7.467 56.987 ;
      VIA 7.422 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 56.413 7.467 56.447 ;
      VIA 7.422 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 55.873 7.467 55.907 ;
      VIA 7.422 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 55.333 7.467 55.367 ;
      VIA 7.422 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 54.793 7.467 54.827 ;
      VIA 7.422 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 54.253 7.467 54.287 ;
      VIA 7.422 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 53.713 7.467 53.747 ;
      VIA 7.422 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 53.173 7.467 53.207 ;
      VIA 7.422 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 52.633 7.467 52.667 ;
      VIA 7.422 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 52.093 7.467 52.127 ;
      VIA 7.422 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 51.553 7.467 51.587 ;
      VIA 7.422 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 51.013 7.467 51.047 ;
      VIA 7.422 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 50.473 7.467 50.507 ;
      VIA 7.422 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 49.933 7.467 49.967 ;
      VIA 7.422 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 49.393 7.467 49.427 ;
      VIA 7.422 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 48.853 7.467 48.887 ;
      VIA 7.422 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 48.313 7.467 48.347 ;
      VIA 7.422 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 47.773 7.467 47.807 ;
      VIA 7.422 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 47.233 7.467 47.267 ;
      VIA 7.422 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 46.693 7.467 46.727 ;
      VIA 7.422 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 46.153 7.467 46.187 ;
      VIA 7.422 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 45.613 7.467 45.647 ;
      VIA 7.422 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 45.073 7.467 45.107 ;
      VIA 7.422 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 44.533 7.467 44.567 ;
      VIA 7.422 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 43.993 7.467 44.027 ;
      VIA 7.422 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 43.453 7.467 43.487 ;
      VIA 7.422 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 42.913 7.467 42.947 ;
      VIA 7.422 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 42.373 7.467 42.407 ;
      VIA 7.422 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 41.833 7.467 41.867 ;
      VIA 7.422 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 41.293 7.467 41.327 ;
      VIA 7.422 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 40.753 7.467 40.787 ;
      VIA 7.422 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 40.213 7.467 40.247 ;
      VIA 7.422 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.673 7.467 39.707 ;
      VIA 7.422 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.133 7.467 39.167 ;
      VIA 7.422 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.593 7.467 38.627 ;
      VIA 7.422 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.053 7.467 38.087 ;
      VIA 7.422 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 37.513 7.467 37.547 ;
      VIA 7.422 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.973 7.467 37.007 ;
      VIA 7.422 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.433 7.467 36.467 ;
      VIA 7.422 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.893 7.467 35.927 ;
      VIA 7.422 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.353 7.467 35.387 ;
      VIA 7.422 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.813 7.467 34.847 ;
      VIA 7.422 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.273 7.467 34.307 ;
      VIA 7.422 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.733 7.467 33.767 ;
      VIA 7.422 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.193 7.467 33.227 ;
      VIA 7.422 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.653 7.467 32.687 ;
      VIA 7.422 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.113 7.467 32.147 ;
      VIA 7.422 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.573 7.467 31.607 ;
      VIA 7.422 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.033 7.467 31.067 ;
      VIA 7.422 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 30.493 7.467 30.527 ;
      VIA 7.422 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.953 7.467 29.987 ;
      VIA 7.422 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.413 7.467 29.447 ;
      VIA 7.422 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.873 7.467 28.907 ;
      VIA 7.422 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.333 7.467 28.367 ;
      VIA 7.422 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.793 7.467 27.827 ;
      VIA 7.422 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.253 7.467 27.287 ;
      VIA 7.422 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.713 7.467 26.747 ;
      VIA 7.422 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.173 7.467 26.207 ;
      VIA 7.422 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.633 7.467 25.667 ;
      VIA 7.422 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.093 7.467 25.127 ;
      VIA 7.422 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.553 7.467 24.587 ;
      VIA 7.422 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.013 7.467 24.047 ;
      VIA 7.422 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 23.473 7.467 23.507 ;
      VIA 7.422 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.933 7.467 22.967 ;
      VIA 7.422 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.393 7.467 22.427 ;
      VIA 7.422 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.853 7.467 21.887 ;
      VIA 7.422 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.313 7.467 21.347 ;
      VIA 7.422 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.773 7.467 20.807 ;
      VIA 7.422 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.233 7.467 20.267 ;
      VIA 7.422 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.693 7.467 19.727 ;
      VIA 7.422 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.153 7.467 19.187 ;
      VIA 7.422 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.613 7.467 18.647 ;
      VIA 7.422 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.073 7.467 18.107 ;
      VIA 7.422 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 17.533 7.467 17.567 ;
      VIA 7.422 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.993 7.467 17.027 ;
      VIA 7.422 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.453 7.467 16.487 ;
      VIA 7.422 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.913 7.467 15.947 ;
      VIA 7.422 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.373 7.467 15.407 ;
      VIA 7.422 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.833 7.467 14.867 ;
      VIA 7.422 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.293 7.467 14.327 ;
      VIA 7.422 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.753 7.467 13.787 ;
      VIA 7.422 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.213 7.467 13.247 ;
      VIA 7.422 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.673 7.467 12.707 ;
      VIA 7.422 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.133 7.467 12.167 ;
      VIA 7.422 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.593 7.467 11.627 ;
      VIA 7.422 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.053 7.467 11.087 ;
      VIA 7.422 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 10.513 7.467 10.547 ;
      VIA 7.422 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.973 7.467 10.007 ;
      VIA 7.422 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.433 7.467 9.467 ;
      VIA 7.422 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.893 7.467 8.927 ;
      VIA 7.422 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.353 7.467 8.387 ;
      VIA 7.422 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.813 7.467 7.847 ;
      VIA 7.422 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.273 7.467 7.307 ;
      VIA 7.422 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.733 7.467 6.767 ;
      VIA 7.422 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.193 7.467 6.227 ;
      VIA 7.422 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.653 7.467 5.687 ;
      VIA 7.422 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.113 7.467 5.147 ;
      VIA 7.422 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.573 7.467 4.607 ;
      VIA 7.422 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.033 7.467 4.067 ;
      VIA 7.422 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 3.493 7.467 3.527 ;
      VIA 7.422 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.953 7.467 2.987 ;
      VIA 7.422 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.413 7.467 2.447 ;
      VIA 7.422 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.873 7.467 1.907 ;
      VIA 7.422 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.333 7.467 1.367 ;
      VIA 7.422 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 73.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 73.153 1.563 73.187 ;
      VIA 1.518 73.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 73.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 72.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 72.613 1.563 72.647 ;
      VIA 1.518 72.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 72.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 72.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 72.073 1.563 72.107 ;
      VIA 1.518 72.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 72.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 71.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 71.533 1.563 71.567 ;
      VIA 1.518 71.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 71.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 71.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 70.993 1.563 71.027 ;
      VIA 1.518 71.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 71.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 70.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 70.453 1.563 70.487 ;
      VIA 1.518 70.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 70.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 69.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 69.913 1.563 69.947 ;
      VIA 1.518 69.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 69.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 69.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 69.373 1.563 69.407 ;
      VIA 1.518 69.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 69.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 68.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 68.833 1.563 68.867 ;
      VIA 1.518 68.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 68.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 68.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 68.293 1.563 68.327 ;
      VIA 1.518 68.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 68.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 67.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 67.753 1.563 67.787 ;
      VIA 1.518 67.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 67.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 67.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 67.213 1.563 67.247 ;
      VIA 1.518 67.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 67.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 66.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 66.673 1.563 66.707 ;
      VIA 1.518 66.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 66.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 66.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 66.133 1.563 66.167 ;
      VIA 1.518 66.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 66.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 65.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 65.593 1.563 65.627 ;
      VIA 1.518 65.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 65.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 65.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 65.053 1.563 65.087 ;
      VIA 1.518 65.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 65.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 64.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 64.513 1.563 64.547 ;
      VIA 1.518 64.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 64.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 63.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 63.973 1.563 64.007 ;
      VIA 1.518 63.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 63.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 63.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 63.433 1.563 63.467 ;
      VIA 1.518 63.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 63.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 62.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 62.893 1.563 62.927 ;
      VIA 1.518 62.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 62.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 62.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 62.353 1.563 62.387 ;
      VIA 1.518 62.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 62.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 61.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 61.813 1.563 61.847 ;
      VIA 1.518 61.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 61.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 61.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 61.273 1.563 61.307 ;
      VIA 1.518 61.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 61.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 60.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 60.733 1.563 60.767 ;
      VIA 1.518 60.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 60.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 60.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 60.193 1.563 60.227 ;
      VIA 1.518 60.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 60.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 59.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 59.653 1.563 59.687 ;
      VIA 1.518 59.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 59.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 59.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 59.113 1.563 59.147 ;
      VIA 1.518 59.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 59.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 58.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 58.573 1.563 58.607 ;
      VIA 1.518 58.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 58.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 58.033 1.563 58.067 ;
      VIA 1.518 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 57.493 1.563 57.527 ;
      VIA 1.518 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 56.953 1.563 56.987 ;
      VIA 1.518 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 56.413 1.563 56.447 ;
      VIA 1.518 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 55.873 1.563 55.907 ;
      VIA 1.518 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 55.333 1.563 55.367 ;
      VIA 1.518 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 54.793 1.563 54.827 ;
      VIA 1.518 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 54.253 1.563 54.287 ;
      VIA 1.518 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 53.713 1.563 53.747 ;
      VIA 1.518 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 53.173 1.563 53.207 ;
      VIA 1.518 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 52.633 1.563 52.667 ;
      VIA 1.518 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 52.093 1.563 52.127 ;
      VIA 1.518 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 51.553 1.563 51.587 ;
      VIA 1.518 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 51.013 1.563 51.047 ;
      VIA 1.518 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 50.473 1.563 50.507 ;
      VIA 1.518 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 49.933 1.563 49.967 ;
      VIA 1.518 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 49.393 1.563 49.427 ;
      VIA 1.518 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 48.853 1.563 48.887 ;
      VIA 1.518 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 48.313 1.563 48.347 ;
      VIA 1.518 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 47.773 1.563 47.807 ;
      VIA 1.518 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 47.233 1.563 47.267 ;
      VIA 1.518 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 46.693 1.563 46.727 ;
      VIA 1.518 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 46.153 1.563 46.187 ;
      VIA 1.518 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 45.613 1.563 45.647 ;
      VIA 1.518 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 45.073 1.563 45.107 ;
      VIA 1.518 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 44.533 1.563 44.567 ;
      VIA 1.518 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 43.993 1.563 44.027 ;
      VIA 1.518 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 43.453 1.563 43.487 ;
      VIA 1.518 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 42.913 1.563 42.947 ;
      VIA 1.518 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 42.373 1.563 42.407 ;
      VIA 1.518 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 41.833 1.563 41.867 ;
      VIA 1.518 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 41.293 1.563 41.327 ;
      VIA 1.518 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 40.753 1.563 40.787 ;
      VIA 1.518 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 40.213 1.563 40.247 ;
      VIA 1.518 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.673 1.563 39.707 ;
      VIA 1.518 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.133 1.563 39.167 ;
      VIA 1.518 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.593 1.563 38.627 ;
      VIA 1.518 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.053 1.563 38.087 ;
      VIA 1.518 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 37.513 1.563 37.547 ;
      VIA 1.518 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.973 1.563 37.007 ;
      VIA 1.518 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.433 1.563 36.467 ;
      VIA 1.518 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.893 1.563 35.927 ;
      VIA 1.518 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.353 1.563 35.387 ;
      VIA 1.518 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.813 1.563 34.847 ;
      VIA 1.518 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.273 1.563 34.307 ;
      VIA 1.518 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.733 1.563 33.767 ;
      VIA 1.518 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.193 1.563 33.227 ;
      VIA 1.518 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.653 1.563 32.687 ;
      VIA 1.518 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.113 1.563 32.147 ;
      VIA 1.518 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.573 1.563 31.607 ;
      VIA 1.518 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.033 1.563 31.067 ;
      VIA 1.518 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 30.493 1.563 30.527 ;
      VIA 1.518 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.953 1.563 29.987 ;
      VIA 1.518 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.413 1.563 29.447 ;
      VIA 1.518 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.873 1.563 28.907 ;
      VIA 1.518 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.333 1.563 28.367 ;
      VIA 1.518 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.793 1.563 27.827 ;
      VIA 1.518 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.253 1.563 27.287 ;
      VIA 1.518 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.713 1.563 26.747 ;
      VIA 1.518 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.173 1.563 26.207 ;
      VIA 1.518 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.633 1.563 25.667 ;
      VIA 1.518 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.093 1.563 25.127 ;
      VIA 1.518 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.553 1.563 24.587 ;
      VIA 1.518 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.013 1.563 24.047 ;
      VIA 1.518 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 23.473 1.563 23.507 ;
      VIA 1.518 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.933 1.563 22.967 ;
      VIA 1.518 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.393 1.563 22.427 ;
      VIA 1.518 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.853 1.563 21.887 ;
      VIA 1.518 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.313 1.563 21.347 ;
      VIA 1.518 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.773 1.563 20.807 ;
      VIA 1.518 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.233 1.563 20.267 ;
      VIA 1.518 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.693 1.563 19.727 ;
      VIA 1.518 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.153 1.563 19.187 ;
      VIA 1.518 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.613 1.563 18.647 ;
      VIA 1.518 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.073 1.563 18.107 ;
      VIA 1.518 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 17.533 1.563 17.567 ;
      VIA 1.518 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.993 1.563 17.027 ;
      VIA 1.518 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.453 1.563 16.487 ;
      VIA 1.518 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.913 1.563 15.947 ;
      VIA 1.518 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.373 1.563 15.407 ;
      VIA 1.518 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.833 1.563 14.867 ;
      VIA 1.518 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.293 1.563 14.327 ;
      VIA 1.518 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.753 1.563 13.787 ;
      VIA 1.518 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.213 1.563 13.247 ;
      VIA 1.518 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.673 1.563 12.707 ;
      VIA 1.518 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.133 1.563 12.167 ;
      VIA 1.518 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.593 1.563 11.627 ;
      VIA 1.518 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.053 1.563 11.087 ;
      VIA 1.518 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 10.513 1.563 10.547 ;
      VIA 1.518 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.973 1.563 10.007 ;
      VIA 1.518 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.433 1.563 9.467 ;
      VIA 1.518 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.893 1.563 8.927 ;
      VIA 1.518 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.353 1.563 8.387 ;
      VIA 1.518 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.813 1.563 7.847 ;
      VIA 1.518 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.273 1.563 7.307 ;
      VIA 1.518 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.733 1.563 6.767 ;
      VIA 1.518 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.193 1.563 6.227 ;
      VIA 1.518 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.653 1.563 5.687 ;
      VIA 1.518 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.113 1.563 5.147 ;
      VIA 1.518 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 37.341 73.17 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 72.63 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 72.09 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 71.55 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 71.01 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 70.47 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 69.93 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 69.39 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 68.85 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 68.31 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 67.77 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 67.23 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 66.69 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 66.15 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 65.61 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 65.07 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 64.53 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 63.99 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 63.45 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 62.91 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 62.37 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 61.83 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 61.29 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 60.75 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 60.21 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 59.67 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 59.13 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 58.59 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 58.05 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 57.51 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 56.97 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 56.43 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 55.89 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 55.35 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 54.81 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 54.27 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 53.73 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 53.19 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 52.65 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 52.11 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 51.57 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 51.03 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 50.49 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 49.95 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 49.41 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 48.87 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 48.33 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 47.79 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 47.25 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 46.71 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 46.17 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 45.63 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 45.09 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 44.55 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 44.01 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 43.47 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 42.93 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 42.39 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 41.85 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 41.31 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 40.77 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 40.23 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 39.69 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 39.15 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 38.61 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 38.07 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 37.53 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 36.99 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 36.45 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 35.91 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 35.37 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 34.83 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 34.29 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 33.75 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 33.21 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 32.67 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 32.13 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 31.59 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 31.05 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 30.51 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 29.97 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 29.43 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 28.89 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 28.35 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 27.81 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 27.27 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 26.73 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 26.19 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 25.65 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 25.11 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 24.57 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 24.03 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 23.49 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 22.95 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 22.41 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 21.87 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 21.33 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 20.79 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 20.25 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 19.71 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 19.17 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 18.63 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 18.09 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 17.55 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 17.01 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 16.47 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 15.93 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 15.39 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 14.85 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 14.31 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 13.77 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 13.23 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 12.69 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 12.15 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 11.61 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 11.07 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 10.53 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 9.99 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 9.45 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 8.91 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 8.37 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 7.83 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 7.29 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 6.75 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 6.21 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 5.67 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 5.13 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 4.59 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 4.05 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 3.51 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 2.97 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 2.43 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 1.89 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 1.35 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.266 67.449 72.234 67.737 ;
        RECT  1.266 61.449 72.234 61.737 ;
        RECT  1.266 55.449 72.234 55.737 ;
        RECT  1.266 49.449 72.234 49.737 ;
        RECT  1.266 43.449 72.234 43.737 ;
        RECT  1.266 37.449 72.234 37.737 ;
        RECT  1.266 31.449 72.234 31.737 ;
        RECT  1.266 25.449 72.234 25.737 ;
        RECT  1.266 19.449 72.234 19.737 ;
        RECT  1.266 13.449 72.234 13.737 ;
        RECT  1.266 7.449 72.234 7.737 ;
        RECT  1.266 1.449 72.234 1.737 ;
      LAYER M5 ;
        RECT  72.114 1.057 72.234 73.463 ;
        RECT  66.21 1.057 66.33 73.463 ;
        RECT  60.306 1.057 60.426 73.463 ;
        RECT  54.402 1.057 54.522 73.463 ;
        RECT  48.498 1.057 48.618 73.463 ;
        RECT  42.594 1.057 42.714 73.463 ;
        RECT  36.69 1.057 36.81 73.463 ;
        RECT  30.786 1.057 30.906 73.463 ;
        RECT  24.882 1.057 25.002 73.463 ;
        RECT  18.978 1.057 19.098 73.463 ;
        RECT  13.074 1.057 13.194 73.463 ;
        RECT  7.17 1.057 7.29 73.463 ;
        RECT  1.266 1.057 1.386 73.463 ;
      LAYER M2 ;
        RECT  1.026 73.431 73.656 73.449 ;
        RECT  1.026 72.891 73.656 72.909 ;
        RECT  1.026 72.351 73.656 72.369 ;
        RECT  1.026 71.811 73.656 71.829 ;
        RECT  1.026 71.271 73.656 71.289 ;
        RECT  1.026 70.731 73.656 70.749 ;
        RECT  1.026 70.191 73.656 70.209 ;
        RECT  1.026 69.651 73.656 69.669 ;
        RECT  1.026 69.111 73.656 69.129 ;
        RECT  1.026 68.571 73.656 68.589 ;
        RECT  1.026 68.031 73.656 68.049 ;
        RECT  1.026 67.491 73.656 67.509 ;
        RECT  1.026 66.951 73.656 66.969 ;
        RECT  1.026 66.411 73.656 66.429 ;
        RECT  1.026 65.871 73.656 65.889 ;
        RECT  1.026 65.331 73.656 65.349 ;
        RECT  1.026 64.791 73.656 64.809 ;
        RECT  1.026 64.251 73.656 64.269 ;
        RECT  1.026 63.711 73.656 63.729 ;
        RECT  1.026 63.171 73.656 63.189 ;
        RECT  1.026 62.631 73.656 62.649 ;
        RECT  1.026 62.091 73.656 62.109 ;
        RECT  1.026 61.551 73.656 61.569 ;
        RECT  1.026 61.011 73.656 61.029 ;
        RECT  1.026 60.471 73.656 60.489 ;
        RECT  1.026 59.931 73.656 59.949 ;
        RECT  1.026 59.391 73.656 59.409 ;
        RECT  1.026 58.851 73.656 58.869 ;
        RECT  1.026 58.311 73.656 58.329 ;
        RECT  1.026 57.771 73.656 57.789 ;
        RECT  1.026 57.231 73.656 57.249 ;
        RECT  1.026 56.691 73.656 56.709 ;
        RECT  1.026 56.151 73.656 56.169 ;
        RECT  1.026 55.611 73.656 55.629 ;
        RECT  1.026 55.071 73.656 55.089 ;
        RECT  1.026 54.531 73.656 54.549 ;
        RECT  1.026 53.991 73.656 54.009 ;
        RECT  1.026 53.451 73.656 53.469 ;
        RECT  1.026 52.911 73.656 52.929 ;
        RECT  1.026 52.371 73.656 52.389 ;
        RECT  1.026 51.831 73.656 51.849 ;
        RECT  1.026 51.291 73.656 51.309 ;
        RECT  1.026 50.751 73.656 50.769 ;
        RECT  1.026 50.211 73.656 50.229 ;
        RECT  1.026 49.671 73.656 49.689 ;
        RECT  1.026 49.131 73.656 49.149 ;
        RECT  1.026 48.591 73.656 48.609 ;
        RECT  1.026 48.051 73.656 48.069 ;
        RECT  1.026 47.511 73.656 47.529 ;
        RECT  1.026 46.971 73.656 46.989 ;
        RECT  1.026 46.431 73.656 46.449 ;
        RECT  1.026 45.891 73.656 45.909 ;
        RECT  1.026 45.351 73.656 45.369 ;
        RECT  1.026 44.811 73.656 44.829 ;
        RECT  1.026 44.271 73.656 44.289 ;
        RECT  1.026 43.731 73.656 43.749 ;
        RECT  1.026 43.191 73.656 43.209 ;
        RECT  1.026 42.651 73.656 42.669 ;
        RECT  1.026 42.111 73.656 42.129 ;
        RECT  1.026 41.571 73.656 41.589 ;
        RECT  1.026 41.031 73.656 41.049 ;
        RECT  1.026 40.491 73.656 40.509 ;
        RECT  1.026 39.951 73.656 39.969 ;
        RECT  1.026 39.411 73.656 39.429 ;
        RECT  1.026 38.871 73.656 38.889 ;
        RECT  1.026 38.331 73.656 38.349 ;
        RECT  1.026 37.791 73.656 37.809 ;
        RECT  1.026 37.251 73.656 37.269 ;
        RECT  1.026 36.711 73.656 36.729 ;
        RECT  1.026 36.171 73.656 36.189 ;
        RECT  1.026 35.631 73.656 35.649 ;
        RECT  1.026 35.091 73.656 35.109 ;
        RECT  1.026 34.551 73.656 34.569 ;
        RECT  1.026 34.011 73.656 34.029 ;
        RECT  1.026 33.471 73.656 33.489 ;
        RECT  1.026 32.931 73.656 32.949 ;
        RECT  1.026 32.391 73.656 32.409 ;
        RECT  1.026 31.851 73.656 31.869 ;
        RECT  1.026 31.311 73.656 31.329 ;
        RECT  1.026 30.771 73.656 30.789 ;
        RECT  1.026 30.231 73.656 30.249 ;
        RECT  1.026 29.691 73.656 29.709 ;
        RECT  1.026 29.151 73.656 29.169 ;
        RECT  1.026 28.611 73.656 28.629 ;
        RECT  1.026 28.071 73.656 28.089 ;
        RECT  1.026 27.531 73.656 27.549 ;
        RECT  1.026 26.991 73.656 27.009 ;
        RECT  1.026 26.451 73.656 26.469 ;
        RECT  1.026 25.911 73.656 25.929 ;
        RECT  1.026 25.371 73.656 25.389 ;
        RECT  1.026 24.831 73.656 24.849 ;
        RECT  1.026 24.291 73.656 24.309 ;
        RECT  1.026 23.751 73.656 23.769 ;
        RECT  1.026 23.211 73.656 23.229 ;
        RECT  1.026 22.671 73.656 22.689 ;
        RECT  1.026 22.131 73.656 22.149 ;
        RECT  1.026 21.591 73.656 21.609 ;
        RECT  1.026 21.051 73.656 21.069 ;
        RECT  1.026 20.511 73.656 20.529 ;
        RECT  1.026 19.971 73.656 19.989 ;
        RECT  1.026 19.431 73.656 19.449 ;
        RECT  1.026 18.891 73.656 18.909 ;
        RECT  1.026 18.351 73.656 18.369 ;
        RECT  1.026 17.811 73.656 17.829 ;
        RECT  1.026 17.271 73.656 17.289 ;
        RECT  1.026 16.731 73.656 16.749 ;
        RECT  1.026 16.191 73.656 16.209 ;
        RECT  1.026 15.651 73.656 15.669 ;
        RECT  1.026 15.111 73.656 15.129 ;
        RECT  1.026 14.571 73.656 14.589 ;
        RECT  1.026 14.031 73.656 14.049 ;
        RECT  1.026 13.491 73.656 13.509 ;
        RECT  1.026 12.951 73.656 12.969 ;
        RECT  1.026 12.411 73.656 12.429 ;
        RECT  1.026 11.871 73.656 11.889 ;
        RECT  1.026 11.331 73.656 11.349 ;
        RECT  1.026 10.791 73.656 10.809 ;
        RECT  1.026 10.251 73.656 10.269 ;
        RECT  1.026 9.711 73.656 9.729 ;
        RECT  1.026 9.171 73.656 9.189 ;
        RECT  1.026 8.631 73.656 8.649 ;
        RECT  1.026 8.091 73.656 8.109 ;
        RECT  1.026 7.551 73.656 7.569 ;
        RECT  1.026 7.011 73.656 7.029 ;
        RECT  1.026 6.471 73.656 6.489 ;
        RECT  1.026 5.931 73.656 5.949 ;
        RECT  1.026 5.391 73.656 5.409 ;
        RECT  1.026 4.851 73.656 4.869 ;
        RECT  1.026 4.311 73.656 4.329 ;
        RECT  1.026 3.771 73.656 3.789 ;
        RECT  1.026 3.231 73.656 3.249 ;
        RECT  1.026 2.691 73.656 2.709 ;
        RECT  1.026 2.151 73.656 2.169 ;
        RECT  1.026 1.611 73.656 1.629 ;
        RECT  1.026 1.071 73.656 1.089 ;
      LAYER M1 ;
        RECT  1.026 73.431 73.656 73.449 ;
        RECT  1.026 72.891 73.656 72.909 ;
        RECT  1.026 72.351 73.656 72.369 ;
        RECT  1.026 71.811 73.656 71.829 ;
        RECT  1.026 71.271 73.656 71.289 ;
        RECT  1.026 70.731 73.656 70.749 ;
        RECT  1.026 70.191 73.656 70.209 ;
        RECT  1.026 69.651 73.656 69.669 ;
        RECT  1.026 69.111 73.656 69.129 ;
        RECT  1.026 68.571 73.656 68.589 ;
        RECT  1.026 68.031 73.656 68.049 ;
        RECT  1.026 67.491 73.656 67.509 ;
        RECT  1.026 66.951 73.656 66.969 ;
        RECT  1.026 66.411 73.656 66.429 ;
        RECT  1.026 65.871 73.656 65.889 ;
        RECT  1.026 65.331 73.656 65.349 ;
        RECT  1.026 64.791 73.656 64.809 ;
        RECT  1.026 64.251 73.656 64.269 ;
        RECT  1.026 63.711 73.656 63.729 ;
        RECT  1.026 63.171 73.656 63.189 ;
        RECT  1.026 62.631 73.656 62.649 ;
        RECT  1.026 62.091 73.656 62.109 ;
        RECT  1.026 61.551 73.656 61.569 ;
        RECT  1.026 61.011 73.656 61.029 ;
        RECT  1.026 60.471 73.656 60.489 ;
        RECT  1.026 59.931 73.656 59.949 ;
        RECT  1.026 59.391 73.656 59.409 ;
        RECT  1.026 58.851 73.656 58.869 ;
        RECT  1.026 58.311 73.656 58.329 ;
        RECT  1.026 57.771 73.656 57.789 ;
        RECT  1.026 57.231 73.656 57.249 ;
        RECT  1.026 56.691 73.656 56.709 ;
        RECT  1.026 56.151 73.656 56.169 ;
        RECT  1.026 55.611 73.656 55.629 ;
        RECT  1.026 55.071 73.656 55.089 ;
        RECT  1.026 54.531 73.656 54.549 ;
        RECT  1.026 53.991 73.656 54.009 ;
        RECT  1.026 53.451 73.656 53.469 ;
        RECT  1.026 52.911 73.656 52.929 ;
        RECT  1.026 52.371 73.656 52.389 ;
        RECT  1.026 51.831 73.656 51.849 ;
        RECT  1.026 51.291 73.656 51.309 ;
        RECT  1.026 50.751 73.656 50.769 ;
        RECT  1.026 50.211 73.656 50.229 ;
        RECT  1.026 49.671 73.656 49.689 ;
        RECT  1.026 49.131 73.656 49.149 ;
        RECT  1.026 48.591 73.656 48.609 ;
        RECT  1.026 48.051 73.656 48.069 ;
        RECT  1.026 47.511 73.656 47.529 ;
        RECT  1.026 46.971 73.656 46.989 ;
        RECT  1.026 46.431 73.656 46.449 ;
        RECT  1.026 45.891 73.656 45.909 ;
        RECT  1.026 45.351 73.656 45.369 ;
        RECT  1.026 44.811 73.656 44.829 ;
        RECT  1.026 44.271 73.656 44.289 ;
        RECT  1.026 43.731 73.656 43.749 ;
        RECT  1.026 43.191 73.656 43.209 ;
        RECT  1.026 42.651 73.656 42.669 ;
        RECT  1.026 42.111 73.656 42.129 ;
        RECT  1.026 41.571 73.656 41.589 ;
        RECT  1.026 41.031 73.656 41.049 ;
        RECT  1.026 40.491 73.656 40.509 ;
        RECT  1.026 39.951 73.656 39.969 ;
        RECT  1.026 39.411 73.656 39.429 ;
        RECT  1.026 38.871 73.656 38.889 ;
        RECT  1.026 38.331 73.656 38.349 ;
        RECT  1.026 37.791 73.656 37.809 ;
        RECT  1.026 37.251 73.656 37.269 ;
        RECT  1.026 36.711 73.656 36.729 ;
        RECT  1.026 36.171 73.656 36.189 ;
        RECT  1.026 35.631 73.656 35.649 ;
        RECT  1.026 35.091 73.656 35.109 ;
        RECT  1.026 34.551 73.656 34.569 ;
        RECT  1.026 34.011 73.656 34.029 ;
        RECT  1.026 33.471 73.656 33.489 ;
        RECT  1.026 32.931 73.656 32.949 ;
        RECT  1.026 32.391 73.656 32.409 ;
        RECT  1.026 31.851 73.656 31.869 ;
        RECT  1.026 31.311 73.656 31.329 ;
        RECT  1.026 30.771 73.656 30.789 ;
        RECT  1.026 30.231 73.656 30.249 ;
        RECT  1.026 29.691 73.656 29.709 ;
        RECT  1.026 29.151 73.656 29.169 ;
        RECT  1.026 28.611 73.656 28.629 ;
        RECT  1.026 28.071 73.656 28.089 ;
        RECT  1.026 27.531 73.656 27.549 ;
        RECT  1.026 26.991 73.656 27.009 ;
        RECT  1.026 26.451 73.656 26.469 ;
        RECT  1.026 25.911 73.656 25.929 ;
        RECT  1.026 25.371 73.656 25.389 ;
        RECT  1.026 24.831 73.656 24.849 ;
        RECT  1.026 24.291 73.656 24.309 ;
        RECT  1.026 23.751 73.656 23.769 ;
        RECT  1.026 23.211 73.656 23.229 ;
        RECT  1.026 22.671 73.656 22.689 ;
        RECT  1.026 22.131 73.656 22.149 ;
        RECT  1.026 21.591 73.656 21.609 ;
        RECT  1.026 21.051 73.656 21.069 ;
        RECT  1.026 20.511 73.656 20.529 ;
        RECT  1.026 19.971 73.656 19.989 ;
        RECT  1.026 19.431 73.656 19.449 ;
        RECT  1.026 18.891 73.656 18.909 ;
        RECT  1.026 18.351 73.656 18.369 ;
        RECT  1.026 17.811 73.656 17.829 ;
        RECT  1.026 17.271 73.656 17.289 ;
        RECT  1.026 16.731 73.656 16.749 ;
        RECT  1.026 16.191 73.656 16.209 ;
        RECT  1.026 15.651 73.656 15.669 ;
        RECT  1.026 15.111 73.656 15.129 ;
        RECT  1.026 14.571 73.656 14.589 ;
        RECT  1.026 14.031 73.656 14.049 ;
        RECT  1.026 13.491 73.656 13.509 ;
        RECT  1.026 12.951 73.656 12.969 ;
        RECT  1.026 12.411 73.656 12.429 ;
        RECT  1.026 11.871 73.656 11.889 ;
        RECT  1.026 11.331 73.656 11.349 ;
        RECT  1.026 10.791 73.656 10.809 ;
        RECT  1.026 10.251 73.656 10.269 ;
        RECT  1.026 9.711 73.656 9.729 ;
        RECT  1.026 9.171 73.656 9.189 ;
        RECT  1.026 8.631 73.656 8.649 ;
        RECT  1.026 8.091 73.656 8.109 ;
        RECT  1.026 7.551 73.656 7.569 ;
        RECT  1.026 7.011 73.656 7.029 ;
        RECT  1.026 6.471 73.656 6.489 ;
        RECT  1.026 5.931 73.656 5.949 ;
        RECT  1.026 5.391 73.656 5.409 ;
        RECT  1.026 4.851 73.656 4.869 ;
        RECT  1.026 4.311 73.656 4.329 ;
        RECT  1.026 3.771 73.656 3.789 ;
        RECT  1.026 3.231 73.656 3.249 ;
        RECT  1.026 2.691 73.656 2.709 ;
        RECT  1.026 2.151 73.656 2.169 ;
        RECT  1.026 1.611 73.656 1.629 ;
        RECT  1.026 1.071 73.656 1.089 ;
      VIA 72.174 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 66.27 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 60.366 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 67.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 61.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 72.174 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 73.423 72.219 73.457 ;
      VIA 72.174 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 72.883 72.219 72.917 ;
      VIA 72.174 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 72.343 72.219 72.377 ;
      VIA 72.174 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 71.803 72.219 71.837 ;
      VIA 72.174 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 71.263 72.219 71.297 ;
      VIA 72.174 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 70.723 72.219 70.757 ;
      VIA 72.174 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 70.183 72.219 70.217 ;
      VIA 72.174 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 69.643 72.219 69.677 ;
      VIA 72.174 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 69.103 72.219 69.137 ;
      VIA 72.174 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 68.563 72.219 68.597 ;
      VIA 72.174 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 68.023 72.219 68.057 ;
      VIA 72.174 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 67.483 72.219 67.517 ;
      VIA 72.174 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 66.943 72.219 66.977 ;
      VIA 72.174 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 66.403 72.219 66.437 ;
      VIA 72.174 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 65.863 72.219 65.897 ;
      VIA 72.174 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 65.323 72.219 65.357 ;
      VIA 72.174 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 64.783 72.219 64.817 ;
      VIA 72.174 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 64.243 72.219 64.277 ;
      VIA 72.174 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 63.703 72.219 63.737 ;
      VIA 72.174 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 63.163 72.219 63.197 ;
      VIA 72.174 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 62.623 72.219 62.657 ;
      VIA 72.174 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 62.083 72.219 62.117 ;
      VIA 72.174 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 61.543 72.219 61.577 ;
      VIA 72.174 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 61.003 72.219 61.037 ;
      VIA 72.174 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 60.463 72.219 60.497 ;
      VIA 72.174 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 59.923 72.219 59.957 ;
      VIA 72.174 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 59.383 72.219 59.417 ;
      VIA 72.174 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 58.843 72.219 58.877 ;
      VIA 72.174 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 58.303 72.219 58.337 ;
      VIA 72.174 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 57.763 72.219 57.797 ;
      VIA 72.174 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 57.223 72.219 57.257 ;
      VIA 72.174 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 56.683 72.219 56.717 ;
      VIA 72.174 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 56.143 72.219 56.177 ;
      VIA 72.174 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 55.603 72.219 55.637 ;
      VIA 72.174 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 55.063 72.219 55.097 ;
      VIA 72.174 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 54.523 72.219 54.557 ;
      VIA 72.174 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 53.983 72.219 54.017 ;
      VIA 72.174 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 53.443 72.219 53.477 ;
      VIA 72.174 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 52.903 72.219 52.937 ;
      VIA 72.174 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 52.363 72.219 52.397 ;
      VIA 72.174 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 51.823 72.219 51.857 ;
      VIA 72.174 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 51.283 72.219 51.317 ;
      VIA 72.174 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 50.743 72.219 50.777 ;
      VIA 72.174 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 50.203 72.219 50.237 ;
      VIA 72.174 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 49.663 72.219 49.697 ;
      VIA 72.174 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 49.123 72.219 49.157 ;
      VIA 72.174 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 48.583 72.219 48.617 ;
      VIA 72.174 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 48.043 72.219 48.077 ;
      VIA 72.174 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 47.503 72.219 47.537 ;
      VIA 72.174 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 46.963 72.219 46.997 ;
      VIA 72.174 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 46.423 72.219 46.457 ;
      VIA 72.174 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 45.883 72.219 45.917 ;
      VIA 72.174 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 45.343 72.219 45.377 ;
      VIA 72.174 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 44.803 72.219 44.837 ;
      VIA 72.174 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 44.263 72.219 44.297 ;
      VIA 72.174 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 43.723 72.219 43.757 ;
      VIA 72.174 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 43.183 72.219 43.217 ;
      VIA 72.174 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 42.643 72.219 42.677 ;
      VIA 72.174 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 42.103 72.219 42.137 ;
      VIA 72.174 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 41.563 72.219 41.597 ;
      VIA 72.174 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 41.023 72.219 41.057 ;
      VIA 72.174 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 40.483 72.219 40.517 ;
      VIA 72.174 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 39.943 72.219 39.977 ;
      VIA 72.174 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 39.403 72.219 39.437 ;
      VIA 72.174 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 38.863 72.219 38.897 ;
      VIA 72.174 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 38.323 72.219 38.357 ;
      VIA 72.174 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 37.783 72.219 37.817 ;
      VIA 72.174 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 37.243 72.219 37.277 ;
      VIA 72.174 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 36.703 72.219 36.737 ;
      VIA 72.174 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 36.163 72.219 36.197 ;
      VIA 72.174 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 35.623 72.219 35.657 ;
      VIA 72.174 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 35.083 72.219 35.117 ;
      VIA 72.174 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 34.543 72.219 34.577 ;
      VIA 72.174 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 34.003 72.219 34.037 ;
      VIA 72.174 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 33.463 72.219 33.497 ;
      VIA 72.174 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 32.923 72.219 32.957 ;
      VIA 72.174 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 32.383 72.219 32.417 ;
      VIA 72.174 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 31.843 72.219 31.877 ;
      VIA 72.174 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 31.303 72.219 31.337 ;
      VIA 72.174 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 30.763 72.219 30.797 ;
      VIA 72.174 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 30.223 72.219 30.257 ;
      VIA 72.174 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 29.683 72.219 29.717 ;
      VIA 72.174 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 29.143 72.219 29.177 ;
      VIA 72.174 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 28.603 72.219 28.637 ;
      VIA 72.174 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 28.063 72.219 28.097 ;
      VIA 72.174 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 27.523 72.219 27.557 ;
      VIA 72.174 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 26.983 72.219 27.017 ;
      VIA 72.174 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 26.443 72.219 26.477 ;
      VIA 72.174 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 25.903 72.219 25.937 ;
      VIA 72.174 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 25.363 72.219 25.397 ;
      VIA 72.174 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 24.823 72.219 24.857 ;
      VIA 72.174 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 24.283 72.219 24.317 ;
      VIA 72.174 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 23.743 72.219 23.777 ;
      VIA 72.174 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 23.203 72.219 23.237 ;
      VIA 72.174 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 22.663 72.219 22.697 ;
      VIA 72.174 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 22.123 72.219 22.157 ;
      VIA 72.174 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 21.583 72.219 21.617 ;
      VIA 72.174 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 21.043 72.219 21.077 ;
      VIA 72.174 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 20.503 72.219 20.537 ;
      VIA 72.174 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 19.963 72.219 19.997 ;
      VIA 72.174 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 19.423 72.219 19.457 ;
      VIA 72.174 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 18.883 72.219 18.917 ;
      VIA 72.174 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 18.343 72.219 18.377 ;
      VIA 72.174 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 17.803 72.219 17.837 ;
      VIA 72.174 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 17.263 72.219 17.297 ;
      VIA 72.174 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 16.723 72.219 16.757 ;
      VIA 72.174 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 16.183 72.219 16.217 ;
      VIA 72.174 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 15.643 72.219 15.677 ;
      VIA 72.174 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 15.103 72.219 15.137 ;
      VIA 72.174 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 14.563 72.219 14.597 ;
      VIA 72.174 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 14.023 72.219 14.057 ;
      VIA 72.174 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 13.483 72.219 13.517 ;
      VIA 72.174 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 12.943 72.219 12.977 ;
      VIA 72.174 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 12.403 72.219 12.437 ;
      VIA 72.174 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 11.863 72.219 11.897 ;
      VIA 72.174 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 11.323 72.219 11.357 ;
      VIA 72.174 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 10.783 72.219 10.817 ;
      VIA 72.174 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 10.243 72.219 10.277 ;
      VIA 72.174 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 9.703 72.219 9.737 ;
      VIA 72.174 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 9.163 72.219 9.197 ;
      VIA 72.174 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 8.623 72.219 8.657 ;
      VIA 72.174 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 8.083 72.219 8.117 ;
      VIA 72.174 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 7.543 72.219 7.577 ;
      VIA 72.174 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 7.003 72.219 7.037 ;
      VIA 72.174 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 6.463 72.219 6.497 ;
      VIA 72.174 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 5.923 72.219 5.957 ;
      VIA 72.174 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 5.383 72.219 5.417 ;
      VIA 72.174 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 4.843 72.219 4.877 ;
      VIA 72.174 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 4.303 72.219 4.337 ;
      VIA 72.174 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 3.763 72.219 3.797 ;
      VIA 72.174 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 3.223 72.219 3.257 ;
      VIA 72.174 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 2.683 72.219 2.717 ;
      VIA 72.174 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 2.143 72.219 2.177 ;
      VIA 72.174 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 1.603 72.219 1.637 ;
      VIA 72.174 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 72.174 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  72.129 1.063 72.219 1.097 ;
      VIA 72.174 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 72.174 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 73.423 66.315 73.457 ;
      VIA 66.27 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 72.883 66.315 72.917 ;
      VIA 66.27 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 72.343 66.315 72.377 ;
      VIA 66.27 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 71.803 66.315 71.837 ;
      VIA 66.27 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 71.263 66.315 71.297 ;
      VIA 66.27 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 70.723 66.315 70.757 ;
      VIA 66.27 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 70.183 66.315 70.217 ;
      VIA 66.27 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 69.643 66.315 69.677 ;
      VIA 66.27 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 69.103 66.315 69.137 ;
      VIA 66.27 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 68.563 66.315 68.597 ;
      VIA 66.27 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 68.023 66.315 68.057 ;
      VIA 66.27 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 67.483 66.315 67.517 ;
      VIA 66.27 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 66.943 66.315 66.977 ;
      VIA 66.27 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 66.403 66.315 66.437 ;
      VIA 66.27 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 65.863 66.315 65.897 ;
      VIA 66.27 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 65.323 66.315 65.357 ;
      VIA 66.27 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 64.783 66.315 64.817 ;
      VIA 66.27 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 64.243 66.315 64.277 ;
      VIA 66.27 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 63.703 66.315 63.737 ;
      VIA 66.27 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 63.163 66.315 63.197 ;
      VIA 66.27 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 62.623 66.315 62.657 ;
      VIA 66.27 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 62.083 66.315 62.117 ;
      VIA 66.27 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 61.543 66.315 61.577 ;
      VIA 66.27 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 61.003 66.315 61.037 ;
      VIA 66.27 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 60.463 66.315 60.497 ;
      VIA 66.27 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 59.923 66.315 59.957 ;
      VIA 66.27 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 59.383 66.315 59.417 ;
      VIA 66.27 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 58.843 66.315 58.877 ;
      VIA 66.27 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 58.303 66.315 58.337 ;
      VIA 66.27 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 57.763 66.315 57.797 ;
      VIA 66.27 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 57.223 66.315 57.257 ;
      VIA 66.27 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 56.683 66.315 56.717 ;
      VIA 66.27 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 56.143 66.315 56.177 ;
      VIA 66.27 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 55.603 66.315 55.637 ;
      VIA 66.27 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 55.063 66.315 55.097 ;
      VIA 66.27 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 54.523 66.315 54.557 ;
      VIA 66.27 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 53.983 66.315 54.017 ;
      VIA 66.27 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 53.443 66.315 53.477 ;
      VIA 66.27 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 52.903 66.315 52.937 ;
      VIA 66.27 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 52.363 66.315 52.397 ;
      VIA 66.27 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 51.823 66.315 51.857 ;
      VIA 66.27 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 51.283 66.315 51.317 ;
      VIA 66.27 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 50.743 66.315 50.777 ;
      VIA 66.27 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 50.203 66.315 50.237 ;
      VIA 66.27 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 49.663 66.315 49.697 ;
      VIA 66.27 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 49.123 66.315 49.157 ;
      VIA 66.27 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 48.583 66.315 48.617 ;
      VIA 66.27 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 48.043 66.315 48.077 ;
      VIA 66.27 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 47.503 66.315 47.537 ;
      VIA 66.27 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 46.963 66.315 46.997 ;
      VIA 66.27 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 46.423 66.315 46.457 ;
      VIA 66.27 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 45.883 66.315 45.917 ;
      VIA 66.27 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 45.343 66.315 45.377 ;
      VIA 66.27 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 44.803 66.315 44.837 ;
      VIA 66.27 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 44.263 66.315 44.297 ;
      VIA 66.27 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 43.723 66.315 43.757 ;
      VIA 66.27 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 43.183 66.315 43.217 ;
      VIA 66.27 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 42.643 66.315 42.677 ;
      VIA 66.27 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 42.103 66.315 42.137 ;
      VIA 66.27 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 41.563 66.315 41.597 ;
      VIA 66.27 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 41.023 66.315 41.057 ;
      VIA 66.27 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 40.483 66.315 40.517 ;
      VIA 66.27 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 39.943 66.315 39.977 ;
      VIA 66.27 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 39.403 66.315 39.437 ;
      VIA 66.27 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 38.863 66.315 38.897 ;
      VIA 66.27 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 38.323 66.315 38.357 ;
      VIA 66.27 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 37.783 66.315 37.817 ;
      VIA 66.27 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 37.243 66.315 37.277 ;
      VIA 66.27 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 36.703 66.315 36.737 ;
      VIA 66.27 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 36.163 66.315 36.197 ;
      VIA 66.27 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 35.623 66.315 35.657 ;
      VIA 66.27 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 35.083 66.315 35.117 ;
      VIA 66.27 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 34.543 66.315 34.577 ;
      VIA 66.27 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 34.003 66.315 34.037 ;
      VIA 66.27 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 33.463 66.315 33.497 ;
      VIA 66.27 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 32.923 66.315 32.957 ;
      VIA 66.27 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 32.383 66.315 32.417 ;
      VIA 66.27 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 31.843 66.315 31.877 ;
      VIA 66.27 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 31.303 66.315 31.337 ;
      VIA 66.27 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 30.763 66.315 30.797 ;
      VIA 66.27 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 30.223 66.315 30.257 ;
      VIA 66.27 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 29.683 66.315 29.717 ;
      VIA 66.27 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 29.143 66.315 29.177 ;
      VIA 66.27 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 28.603 66.315 28.637 ;
      VIA 66.27 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 28.063 66.315 28.097 ;
      VIA 66.27 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 27.523 66.315 27.557 ;
      VIA 66.27 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 26.983 66.315 27.017 ;
      VIA 66.27 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 26.443 66.315 26.477 ;
      VIA 66.27 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 25.903 66.315 25.937 ;
      VIA 66.27 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 25.363 66.315 25.397 ;
      VIA 66.27 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 24.823 66.315 24.857 ;
      VIA 66.27 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 24.283 66.315 24.317 ;
      VIA 66.27 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 23.743 66.315 23.777 ;
      VIA 66.27 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 23.203 66.315 23.237 ;
      VIA 66.27 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 22.663 66.315 22.697 ;
      VIA 66.27 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 22.123 66.315 22.157 ;
      VIA 66.27 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 21.583 66.315 21.617 ;
      VIA 66.27 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 21.043 66.315 21.077 ;
      VIA 66.27 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 20.503 66.315 20.537 ;
      VIA 66.27 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 19.963 66.315 19.997 ;
      VIA 66.27 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 19.423 66.315 19.457 ;
      VIA 66.27 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 18.883 66.315 18.917 ;
      VIA 66.27 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 18.343 66.315 18.377 ;
      VIA 66.27 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 17.803 66.315 17.837 ;
      VIA 66.27 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 17.263 66.315 17.297 ;
      VIA 66.27 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 16.723 66.315 16.757 ;
      VIA 66.27 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 16.183 66.315 16.217 ;
      VIA 66.27 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 15.643 66.315 15.677 ;
      VIA 66.27 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 15.103 66.315 15.137 ;
      VIA 66.27 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 14.563 66.315 14.597 ;
      VIA 66.27 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 14.023 66.315 14.057 ;
      VIA 66.27 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 13.483 66.315 13.517 ;
      VIA 66.27 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 12.943 66.315 12.977 ;
      VIA 66.27 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 12.403 66.315 12.437 ;
      VIA 66.27 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 11.863 66.315 11.897 ;
      VIA 66.27 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 11.323 66.315 11.357 ;
      VIA 66.27 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 10.783 66.315 10.817 ;
      VIA 66.27 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 10.243 66.315 10.277 ;
      VIA 66.27 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 9.703 66.315 9.737 ;
      VIA 66.27 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 9.163 66.315 9.197 ;
      VIA 66.27 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 8.623 66.315 8.657 ;
      VIA 66.27 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 8.083 66.315 8.117 ;
      VIA 66.27 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 7.543 66.315 7.577 ;
      VIA 66.27 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 7.003 66.315 7.037 ;
      VIA 66.27 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 6.463 66.315 6.497 ;
      VIA 66.27 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 5.923 66.315 5.957 ;
      VIA 66.27 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 5.383 66.315 5.417 ;
      VIA 66.27 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 4.843 66.315 4.877 ;
      VIA 66.27 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 4.303 66.315 4.337 ;
      VIA 66.27 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 3.763 66.315 3.797 ;
      VIA 66.27 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 3.223 66.315 3.257 ;
      VIA 66.27 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 2.683 66.315 2.717 ;
      VIA 66.27 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 2.143 66.315 2.177 ;
      VIA 66.27 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 1.603 66.315 1.637 ;
      VIA 66.27 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 66.27 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  66.225 1.063 66.315 1.097 ;
      VIA 66.27 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 66.27 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 73.423 60.411 73.457 ;
      VIA 60.366 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 72.883 60.411 72.917 ;
      VIA 60.366 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 72.343 60.411 72.377 ;
      VIA 60.366 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 71.803 60.411 71.837 ;
      VIA 60.366 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 71.263 60.411 71.297 ;
      VIA 60.366 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 70.723 60.411 70.757 ;
      VIA 60.366 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 70.183 60.411 70.217 ;
      VIA 60.366 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 69.643 60.411 69.677 ;
      VIA 60.366 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 69.103 60.411 69.137 ;
      VIA 60.366 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 68.563 60.411 68.597 ;
      VIA 60.366 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 68.023 60.411 68.057 ;
      VIA 60.366 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 67.483 60.411 67.517 ;
      VIA 60.366 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 66.943 60.411 66.977 ;
      VIA 60.366 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 66.403 60.411 66.437 ;
      VIA 60.366 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 65.863 60.411 65.897 ;
      VIA 60.366 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 65.323 60.411 65.357 ;
      VIA 60.366 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 64.783 60.411 64.817 ;
      VIA 60.366 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 64.243 60.411 64.277 ;
      VIA 60.366 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 63.703 60.411 63.737 ;
      VIA 60.366 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 63.163 60.411 63.197 ;
      VIA 60.366 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 62.623 60.411 62.657 ;
      VIA 60.366 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 62.083 60.411 62.117 ;
      VIA 60.366 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 61.543 60.411 61.577 ;
      VIA 60.366 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 61.003 60.411 61.037 ;
      VIA 60.366 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 60.463 60.411 60.497 ;
      VIA 60.366 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 59.923 60.411 59.957 ;
      VIA 60.366 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 59.383 60.411 59.417 ;
      VIA 60.366 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 58.843 60.411 58.877 ;
      VIA 60.366 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 58.303 60.411 58.337 ;
      VIA 60.366 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 57.763 60.411 57.797 ;
      VIA 60.366 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 57.223 60.411 57.257 ;
      VIA 60.366 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 56.683 60.411 56.717 ;
      VIA 60.366 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 56.143 60.411 56.177 ;
      VIA 60.366 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 55.603 60.411 55.637 ;
      VIA 60.366 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 55.063 60.411 55.097 ;
      VIA 60.366 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 54.523 60.411 54.557 ;
      VIA 60.366 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 53.983 60.411 54.017 ;
      VIA 60.366 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 53.443 60.411 53.477 ;
      VIA 60.366 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 52.903 60.411 52.937 ;
      VIA 60.366 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 52.363 60.411 52.397 ;
      VIA 60.366 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 51.823 60.411 51.857 ;
      VIA 60.366 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 51.283 60.411 51.317 ;
      VIA 60.366 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 50.743 60.411 50.777 ;
      VIA 60.366 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 50.203 60.411 50.237 ;
      VIA 60.366 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 49.663 60.411 49.697 ;
      VIA 60.366 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 49.123 60.411 49.157 ;
      VIA 60.366 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 48.583 60.411 48.617 ;
      VIA 60.366 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 48.043 60.411 48.077 ;
      VIA 60.366 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 47.503 60.411 47.537 ;
      VIA 60.366 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 46.963 60.411 46.997 ;
      VIA 60.366 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 46.423 60.411 46.457 ;
      VIA 60.366 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 45.883 60.411 45.917 ;
      VIA 60.366 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 45.343 60.411 45.377 ;
      VIA 60.366 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 44.803 60.411 44.837 ;
      VIA 60.366 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 44.263 60.411 44.297 ;
      VIA 60.366 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 43.723 60.411 43.757 ;
      VIA 60.366 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 43.183 60.411 43.217 ;
      VIA 60.366 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 42.643 60.411 42.677 ;
      VIA 60.366 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 42.103 60.411 42.137 ;
      VIA 60.366 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 41.563 60.411 41.597 ;
      VIA 60.366 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 41.023 60.411 41.057 ;
      VIA 60.366 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 40.483 60.411 40.517 ;
      VIA 60.366 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 39.943 60.411 39.977 ;
      VIA 60.366 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 39.403 60.411 39.437 ;
      VIA 60.366 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 38.863 60.411 38.897 ;
      VIA 60.366 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 38.323 60.411 38.357 ;
      VIA 60.366 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 37.783 60.411 37.817 ;
      VIA 60.366 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 37.243 60.411 37.277 ;
      VIA 60.366 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 36.703 60.411 36.737 ;
      VIA 60.366 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 36.163 60.411 36.197 ;
      VIA 60.366 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 35.623 60.411 35.657 ;
      VIA 60.366 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 35.083 60.411 35.117 ;
      VIA 60.366 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 34.543 60.411 34.577 ;
      VIA 60.366 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 34.003 60.411 34.037 ;
      VIA 60.366 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 33.463 60.411 33.497 ;
      VIA 60.366 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 32.923 60.411 32.957 ;
      VIA 60.366 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 32.383 60.411 32.417 ;
      VIA 60.366 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 31.843 60.411 31.877 ;
      VIA 60.366 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 31.303 60.411 31.337 ;
      VIA 60.366 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 30.763 60.411 30.797 ;
      VIA 60.366 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 30.223 60.411 30.257 ;
      VIA 60.366 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 29.683 60.411 29.717 ;
      VIA 60.366 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 29.143 60.411 29.177 ;
      VIA 60.366 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 28.603 60.411 28.637 ;
      VIA 60.366 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 28.063 60.411 28.097 ;
      VIA 60.366 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 27.523 60.411 27.557 ;
      VIA 60.366 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 26.983 60.411 27.017 ;
      VIA 60.366 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 26.443 60.411 26.477 ;
      VIA 60.366 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 25.903 60.411 25.937 ;
      VIA 60.366 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 25.363 60.411 25.397 ;
      VIA 60.366 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 24.823 60.411 24.857 ;
      VIA 60.366 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 24.283 60.411 24.317 ;
      VIA 60.366 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 23.743 60.411 23.777 ;
      VIA 60.366 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 23.203 60.411 23.237 ;
      VIA 60.366 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 22.663 60.411 22.697 ;
      VIA 60.366 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 22.123 60.411 22.157 ;
      VIA 60.366 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 21.583 60.411 21.617 ;
      VIA 60.366 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 21.043 60.411 21.077 ;
      VIA 60.366 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 20.503 60.411 20.537 ;
      VIA 60.366 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 19.963 60.411 19.997 ;
      VIA 60.366 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 19.423 60.411 19.457 ;
      VIA 60.366 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 18.883 60.411 18.917 ;
      VIA 60.366 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 18.343 60.411 18.377 ;
      VIA 60.366 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 17.803 60.411 17.837 ;
      VIA 60.366 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 17.263 60.411 17.297 ;
      VIA 60.366 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 16.723 60.411 16.757 ;
      VIA 60.366 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 16.183 60.411 16.217 ;
      VIA 60.366 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 15.643 60.411 15.677 ;
      VIA 60.366 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 15.103 60.411 15.137 ;
      VIA 60.366 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 14.563 60.411 14.597 ;
      VIA 60.366 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 14.023 60.411 14.057 ;
      VIA 60.366 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 13.483 60.411 13.517 ;
      VIA 60.366 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 12.943 60.411 12.977 ;
      VIA 60.366 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 12.403 60.411 12.437 ;
      VIA 60.366 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 11.863 60.411 11.897 ;
      VIA 60.366 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 11.323 60.411 11.357 ;
      VIA 60.366 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 10.783 60.411 10.817 ;
      VIA 60.366 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 10.243 60.411 10.277 ;
      VIA 60.366 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 9.703 60.411 9.737 ;
      VIA 60.366 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 9.163 60.411 9.197 ;
      VIA 60.366 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 8.623 60.411 8.657 ;
      VIA 60.366 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 8.083 60.411 8.117 ;
      VIA 60.366 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 7.543 60.411 7.577 ;
      VIA 60.366 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 7.003 60.411 7.037 ;
      VIA 60.366 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 6.463 60.411 6.497 ;
      VIA 60.366 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 5.923 60.411 5.957 ;
      VIA 60.366 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 5.383 60.411 5.417 ;
      VIA 60.366 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 4.843 60.411 4.877 ;
      VIA 60.366 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 4.303 60.411 4.337 ;
      VIA 60.366 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 3.763 60.411 3.797 ;
      VIA 60.366 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 3.223 60.411 3.257 ;
      VIA 60.366 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 2.683 60.411 2.717 ;
      VIA 60.366 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 2.143 60.411 2.177 ;
      VIA 60.366 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 1.603 60.411 1.637 ;
      VIA 60.366 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 60.366 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  60.321 1.063 60.411 1.097 ;
      VIA 60.366 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 60.366 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 73.423 54.507 73.457 ;
      VIA 54.462 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 72.883 54.507 72.917 ;
      VIA 54.462 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 72.343 54.507 72.377 ;
      VIA 54.462 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 71.803 54.507 71.837 ;
      VIA 54.462 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 71.263 54.507 71.297 ;
      VIA 54.462 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 70.723 54.507 70.757 ;
      VIA 54.462 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 70.183 54.507 70.217 ;
      VIA 54.462 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 69.643 54.507 69.677 ;
      VIA 54.462 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 69.103 54.507 69.137 ;
      VIA 54.462 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 68.563 54.507 68.597 ;
      VIA 54.462 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 68.023 54.507 68.057 ;
      VIA 54.462 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 67.483 54.507 67.517 ;
      VIA 54.462 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 66.943 54.507 66.977 ;
      VIA 54.462 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 66.403 54.507 66.437 ;
      VIA 54.462 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 65.863 54.507 65.897 ;
      VIA 54.462 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 65.323 54.507 65.357 ;
      VIA 54.462 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 64.783 54.507 64.817 ;
      VIA 54.462 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 64.243 54.507 64.277 ;
      VIA 54.462 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 63.703 54.507 63.737 ;
      VIA 54.462 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 63.163 54.507 63.197 ;
      VIA 54.462 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 62.623 54.507 62.657 ;
      VIA 54.462 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 62.083 54.507 62.117 ;
      VIA 54.462 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 61.543 54.507 61.577 ;
      VIA 54.462 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 61.003 54.507 61.037 ;
      VIA 54.462 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 60.463 54.507 60.497 ;
      VIA 54.462 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 59.923 54.507 59.957 ;
      VIA 54.462 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 59.383 54.507 59.417 ;
      VIA 54.462 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 58.843 54.507 58.877 ;
      VIA 54.462 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 58.303 54.507 58.337 ;
      VIA 54.462 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 57.763 54.507 57.797 ;
      VIA 54.462 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 57.223 54.507 57.257 ;
      VIA 54.462 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 56.683 54.507 56.717 ;
      VIA 54.462 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 56.143 54.507 56.177 ;
      VIA 54.462 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 55.603 54.507 55.637 ;
      VIA 54.462 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 55.063 54.507 55.097 ;
      VIA 54.462 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 54.523 54.507 54.557 ;
      VIA 54.462 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 53.983 54.507 54.017 ;
      VIA 54.462 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 53.443 54.507 53.477 ;
      VIA 54.462 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 52.903 54.507 52.937 ;
      VIA 54.462 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 52.363 54.507 52.397 ;
      VIA 54.462 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 51.823 54.507 51.857 ;
      VIA 54.462 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 51.283 54.507 51.317 ;
      VIA 54.462 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 50.743 54.507 50.777 ;
      VIA 54.462 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 50.203 54.507 50.237 ;
      VIA 54.462 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 49.663 54.507 49.697 ;
      VIA 54.462 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 49.123 54.507 49.157 ;
      VIA 54.462 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 48.583 54.507 48.617 ;
      VIA 54.462 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 48.043 54.507 48.077 ;
      VIA 54.462 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 47.503 54.507 47.537 ;
      VIA 54.462 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 46.963 54.507 46.997 ;
      VIA 54.462 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 46.423 54.507 46.457 ;
      VIA 54.462 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 45.883 54.507 45.917 ;
      VIA 54.462 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 45.343 54.507 45.377 ;
      VIA 54.462 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 44.803 54.507 44.837 ;
      VIA 54.462 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 44.263 54.507 44.297 ;
      VIA 54.462 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 43.723 54.507 43.757 ;
      VIA 54.462 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 43.183 54.507 43.217 ;
      VIA 54.462 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 42.643 54.507 42.677 ;
      VIA 54.462 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 42.103 54.507 42.137 ;
      VIA 54.462 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 41.563 54.507 41.597 ;
      VIA 54.462 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 41.023 54.507 41.057 ;
      VIA 54.462 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 40.483 54.507 40.517 ;
      VIA 54.462 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 39.943 54.507 39.977 ;
      VIA 54.462 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 39.403 54.507 39.437 ;
      VIA 54.462 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 38.863 54.507 38.897 ;
      VIA 54.462 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 38.323 54.507 38.357 ;
      VIA 54.462 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 37.783 54.507 37.817 ;
      VIA 54.462 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 37.243 54.507 37.277 ;
      VIA 54.462 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 36.703 54.507 36.737 ;
      VIA 54.462 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 36.163 54.507 36.197 ;
      VIA 54.462 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 35.623 54.507 35.657 ;
      VIA 54.462 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 35.083 54.507 35.117 ;
      VIA 54.462 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 34.543 54.507 34.577 ;
      VIA 54.462 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 34.003 54.507 34.037 ;
      VIA 54.462 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 33.463 54.507 33.497 ;
      VIA 54.462 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 32.923 54.507 32.957 ;
      VIA 54.462 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 32.383 54.507 32.417 ;
      VIA 54.462 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 31.843 54.507 31.877 ;
      VIA 54.462 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 31.303 54.507 31.337 ;
      VIA 54.462 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 30.763 54.507 30.797 ;
      VIA 54.462 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 30.223 54.507 30.257 ;
      VIA 54.462 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 29.683 54.507 29.717 ;
      VIA 54.462 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 29.143 54.507 29.177 ;
      VIA 54.462 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 28.603 54.507 28.637 ;
      VIA 54.462 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 28.063 54.507 28.097 ;
      VIA 54.462 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 27.523 54.507 27.557 ;
      VIA 54.462 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 26.983 54.507 27.017 ;
      VIA 54.462 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 26.443 54.507 26.477 ;
      VIA 54.462 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 25.903 54.507 25.937 ;
      VIA 54.462 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 25.363 54.507 25.397 ;
      VIA 54.462 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 24.823 54.507 24.857 ;
      VIA 54.462 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 24.283 54.507 24.317 ;
      VIA 54.462 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 23.743 54.507 23.777 ;
      VIA 54.462 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 23.203 54.507 23.237 ;
      VIA 54.462 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 22.663 54.507 22.697 ;
      VIA 54.462 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 22.123 54.507 22.157 ;
      VIA 54.462 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 21.583 54.507 21.617 ;
      VIA 54.462 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 21.043 54.507 21.077 ;
      VIA 54.462 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 20.503 54.507 20.537 ;
      VIA 54.462 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 19.963 54.507 19.997 ;
      VIA 54.462 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 19.423 54.507 19.457 ;
      VIA 54.462 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 18.883 54.507 18.917 ;
      VIA 54.462 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 18.343 54.507 18.377 ;
      VIA 54.462 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 17.803 54.507 17.837 ;
      VIA 54.462 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 17.263 54.507 17.297 ;
      VIA 54.462 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 16.723 54.507 16.757 ;
      VIA 54.462 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 16.183 54.507 16.217 ;
      VIA 54.462 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 15.643 54.507 15.677 ;
      VIA 54.462 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 15.103 54.507 15.137 ;
      VIA 54.462 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 14.563 54.507 14.597 ;
      VIA 54.462 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 14.023 54.507 14.057 ;
      VIA 54.462 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 13.483 54.507 13.517 ;
      VIA 54.462 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 12.943 54.507 12.977 ;
      VIA 54.462 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 12.403 54.507 12.437 ;
      VIA 54.462 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 11.863 54.507 11.897 ;
      VIA 54.462 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 11.323 54.507 11.357 ;
      VIA 54.462 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 10.783 54.507 10.817 ;
      VIA 54.462 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 10.243 54.507 10.277 ;
      VIA 54.462 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 9.703 54.507 9.737 ;
      VIA 54.462 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 9.163 54.507 9.197 ;
      VIA 54.462 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 8.623 54.507 8.657 ;
      VIA 54.462 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 8.083 54.507 8.117 ;
      VIA 54.462 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 7.543 54.507 7.577 ;
      VIA 54.462 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 7.003 54.507 7.037 ;
      VIA 54.462 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 6.463 54.507 6.497 ;
      VIA 54.462 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 5.923 54.507 5.957 ;
      VIA 54.462 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 5.383 54.507 5.417 ;
      VIA 54.462 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 4.843 54.507 4.877 ;
      VIA 54.462 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 4.303 54.507 4.337 ;
      VIA 54.462 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 3.763 54.507 3.797 ;
      VIA 54.462 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 3.223 54.507 3.257 ;
      VIA 54.462 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 2.683 54.507 2.717 ;
      VIA 54.462 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 2.143 54.507 2.177 ;
      VIA 54.462 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 1.603 54.507 1.637 ;
      VIA 54.462 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 1.063 54.507 1.097 ;
      VIA 54.462 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 73.423 48.603 73.457 ;
      VIA 48.558 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 72.883 48.603 72.917 ;
      VIA 48.558 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 72.343 48.603 72.377 ;
      VIA 48.558 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 71.803 48.603 71.837 ;
      VIA 48.558 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 71.263 48.603 71.297 ;
      VIA 48.558 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 70.723 48.603 70.757 ;
      VIA 48.558 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 70.183 48.603 70.217 ;
      VIA 48.558 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 69.643 48.603 69.677 ;
      VIA 48.558 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 69.103 48.603 69.137 ;
      VIA 48.558 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 68.563 48.603 68.597 ;
      VIA 48.558 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 68.023 48.603 68.057 ;
      VIA 48.558 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 67.483 48.603 67.517 ;
      VIA 48.558 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 66.943 48.603 66.977 ;
      VIA 48.558 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 66.403 48.603 66.437 ;
      VIA 48.558 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 65.863 48.603 65.897 ;
      VIA 48.558 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 65.323 48.603 65.357 ;
      VIA 48.558 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 64.783 48.603 64.817 ;
      VIA 48.558 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 64.243 48.603 64.277 ;
      VIA 48.558 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 63.703 48.603 63.737 ;
      VIA 48.558 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 63.163 48.603 63.197 ;
      VIA 48.558 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 62.623 48.603 62.657 ;
      VIA 48.558 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 62.083 48.603 62.117 ;
      VIA 48.558 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 61.543 48.603 61.577 ;
      VIA 48.558 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 61.003 48.603 61.037 ;
      VIA 48.558 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 60.463 48.603 60.497 ;
      VIA 48.558 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 59.923 48.603 59.957 ;
      VIA 48.558 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 59.383 48.603 59.417 ;
      VIA 48.558 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 58.843 48.603 58.877 ;
      VIA 48.558 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 58.303 48.603 58.337 ;
      VIA 48.558 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 57.763 48.603 57.797 ;
      VIA 48.558 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 57.223 48.603 57.257 ;
      VIA 48.558 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 56.683 48.603 56.717 ;
      VIA 48.558 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 56.143 48.603 56.177 ;
      VIA 48.558 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 55.603 48.603 55.637 ;
      VIA 48.558 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 55.063 48.603 55.097 ;
      VIA 48.558 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 54.523 48.603 54.557 ;
      VIA 48.558 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 53.983 48.603 54.017 ;
      VIA 48.558 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 53.443 48.603 53.477 ;
      VIA 48.558 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 52.903 48.603 52.937 ;
      VIA 48.558 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 52.363 48.603 52.397 ;
      VIA 48.558 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 51.823 48.603 51.857 ;
      VIA 48.558 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 51.283 48.603 51.317 ;
      VIA 48.558 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 50.743 48.603 50.777 ;
      VIA 48.558 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 50.203 48.603 50.237 ;
      VIA 48.558 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 49.663 48.603 49.697 ;
      VIA 48.558 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 49.123 48.603 49.157 ;
      VIA 48.558 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 48.583 48.603 48.617 ;
      VIA 48.558 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 48.043 48.603 48.077 ;
      VIA 48.558 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 47.503 48.603 47.537 ;
      VIA 48.558 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 46.963 48.603 46.997 ;
      VIA 48.558 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 46.423 48.603 46.457 ;
      VIA 48.558 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 45.883 48.603 45.917 ;
      VIA 48.558 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 45.343 48.603 45.377 ;
      VIA 48.558 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 44.803 48.603 44.837 ;
      VIA 48.558 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 44.263 48.603 44.297 ;
      VIA 48.558 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 43.723 48.603 43.757 ;
      VIA 48.558 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 43.183 48.603 43.217 ;
      VIA 48.558 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 42.643 48.603 42.677 ;
      VIA 48.558 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 42.103 48.603 42.137 ;
      VIA 48.558 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 41.563 48.603 41.597 ;
      VIA 48.558 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 41.023 48.603 41.057 ;
      VIA 48.558 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 40.483 48.603 40.517 ;
      VIA 48.558 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 39.943 48.603 39.977 ;
      VIA 48.558 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 39.403 48.603 39.437 ;
      VIA 48.558 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 38.863 48.603 38.897 ;
      VIA 48.558 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 38.323 48.603 38.357 ;
      VIA 48.558 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 37.783 48.603 37.817 ;
      VIA 48.558 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 37.243 48.603 37.277 ;
      VIA 48.558 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 36.703 48.603 36.737 ;
      VIA 48.558 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 36.163 48.603 36.197 ;
      VIA 48.558 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 35.623 48.603 35.657 ;
      VIA 48.558 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 35.083 48.603 35.117 ;
      VIA 48.558 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 34.543 48.603 34.577 ;
      VIA 48.558 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 34.003 48.603 34.037 ;
      VIA 48.558 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 33.463 48.603 33.497 ;
      VIA 48.558 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 32.923 48.603 32.957 ;
      VIA 48.558 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 32.383 48.603 32.417 ;
      VIA 48.558 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 31.843 48.603 31.877 ;
      VIA 48.558 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 31.303 48.603 31.337 ;
      VIA 48.558 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 30.763 48.603 30.797 ;
      VIA 48.558 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 30.223 48.603 30.257 ;
      VIA 48.558 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 29.683 48.603 29.717 ;
      VIA 48.558 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 29.143 48.603 29.177 ;
      VIA 48.558 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 28.603 48.603 28.637 ;
      VIA 48.558 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 28.063 48.603 28.097 ;
      VIA 48.558 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 27.523 48.603 27.557 ;
      VIA 48.558 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 26.983 48.603 27.017 ;
      VIA 48.558 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 26.443 48.603 26.477 ;
      VIA 48.558 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 25.903 48.603 25.937 ;
      VIA 48.558 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 25.363 48.603 25.397 ;
      VIA 48.558 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 24.823 48.603 24.857 ;
      VIA 48.558 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 24.283 48.603 24.317 ;
      VIA 48.558 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 23.743 48.603 23.777 ;
      VIA 48.558 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 23.203 48.603 23.237 ;
      VIA 48.558 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 22.663 48.603 22.697 ;
      VIA 48.558 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 22.123 48.603 22.157 ;
      VIA 48.558 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 21.583 48.603 21.617 ;
      VIA 48.558 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 21.043 48.603 21.077 ;
      VIA 48.558 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 20.503 48.603 20.537 ;
      VIA 48.558 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 19.963 48.603 19.997 ;
      VIA 48.558 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 19.423 48.603 19.457 ;
      VIA 48.558 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 18.883 48.603 18.917 ;
      VIA 48.558 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 18.343 48.603 18.377 ;
      VIA 48.558 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 17.803 48.603 17.837 ;
      VIA 48.558 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 17.263 48.603 17.297 ;
      VIA 48.558 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 16.723 48.603 16.757 ;
      VIA 48.558 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 16.183 48.603 16.217 ;
      VIA 48.558 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 15.643 48.603 15.677 ;
      VIA 48.558 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 15.103 48.603 15.137 ;
      VIA 48.558 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 14.563 48.603 14.597 ;
      VIA 48.558 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 14.023 48.603 14.057 ;
      VIA 48.558 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 13.483 48.603 13.517 ;
      VIA 48.558 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 12.943 48.603 12.977 ;
      VIA 48.558 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 12.403 48.603 12.437 ;
      VIA 48.558 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 11.863 48.603 11.897 ;
      VIA 48.558 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 11.323 48.603 11.357 ;
      VIA 48.558 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 10.783 48.603 10.817 ;
      VIA 48.558 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 10.243 48.603 10.277 ;
      VIA 48.558 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 9.703 48.603 9.737 ;
      VIA 48.558 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 9.163 48.603 9.197 ;
      VIA 48.558 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 8.623 48.603 8.657 ;
      VIA 48.558 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 8.083 48.603 8.117 ;
      VIA 48.558 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 7.543 48.603 7.577 ;
      VIA 48.558 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 7.003 48.603 7.037 ;
      VIA 48.558 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 6.463 48.603 6.497 ;
      VIA 48.558 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 5.923 48.603 5.957 ;
      VIA 48.558 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 5.383 48.603 5.417 ;
      VIA 48.558 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 4.843 48.603 4.877 ;
      VIA 48.558 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 4.303 48.603 4.337 ;
      VIA 48.558 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 3.763 48.603 3.797 ;
      VIA 48.558 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 3.223 48.603 3.257 ;
      VIA 48.558 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 2.683 48.603 2.717 ;
      VIA 48.558 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 2.143 48.603 2.177 ;
      VIA 48.558 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 1.603 48.603 1.637 ;
      VIA 48.558 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 1.063 48.603 1.097 ;
      VIA 48.558 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 73.423 42.699 73.457 ;
      VIA 42.654 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 72.883 42.699 72.917 ;
      VIA 42.654 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 72.343 42.699 72.377 ;
      VIA 42.654 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 71.803 42.699 71.837 ;
      VIA 42.654 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 71.263 42.699 71.297 ;
      VIA 42.654 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 70.723 42.699 70.757 ;
      VIA 42.654 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 70.183 42.699 70.217 ;
      VIA 42.654 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 69.643 42.699 69.677 ;
      VIA 42.654 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 69.103 42.699 69.137 ;
      VIA 42.654 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 68.563 42.699 68.597 ;
      VIA 42.654 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 68.023 42.699 68.057 ;
      VIA 42.654 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 67.483 42.699 67.517 ;
      VIA 42.654 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 66.943 42.699 66.977 ;
      VIA 42.654 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 66.403 42.699 66.437 ;
      VIA 42.654 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 65.863 42.699 65.897 ;
      VIA 42.654 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 65.323 42.699 65.357 ;
      VIA 42.654 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 64.783 42.699 64.817 ;
      VIA 42.654 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 64.243 42.699 64.277 ;
      VIA 42.654 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 63.703 42.699 63.737 ;
      VIA 42.654 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 63.163 42.699 63.197 ;
      VIA 42.654 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 62.623 42.699 62.657 ;
      VIA 42.654 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 62.083 42.699 62.117 ;
      VIA 42.654 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 61.543 42.699 61.577 ;
      VIA 42.654 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 61.003 42.699 61.037 ;
      VIA 42.654 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 60.463 42.699 60.497 ;
      VIA 42.654 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 59.923 42.699 59.957 ;
      VIA 42.654 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 59.383 42.699 59.417 ;
      VIA 42.654 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 58.843 42.699 58.877 ;
      VIA 42.654 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 58.303 42.699 58.337 ;
      VIA 42.654 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 57.763 42.699 57.797 ;
      VIA 42.654 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 57.223 42.699 57.257 ;
      VIA 42.654 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 56.683 42.699 56.717 ;
      VIA 42.654 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 56.143 42.699 56.177 ;
      VIA 42.654 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 55.603 42.699 55.637 ;
      VIA 42.654 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 55.063 42.699 55.097 ;
      VIA 42.654 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 54.523 42.699 54.557 ;
      VIA 42.654 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 53.983 42.699 54.017 ;
      VIA 42.654 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 53.443 42.699 53.477 ;
      VIA 42.654 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 52.903 42.699 52.937 ;
      VIA 42.654 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 52.363 42.699 52.397 ;
      VIA 42.654 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 51.823 42.699 51.857 ;
      VIA 42.654 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 51.283 42.699 51.317 ;
      VIA 42.654 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 50.743 42.699 50.777 ;
      VIA 42.654 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 50.203 42.699 50.237 ;
      VIA 42.654 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 49.663 42.699 49.697 ;
      VIA 42.654 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 49.123 42.699 49.157 ;
      VIA 42.654 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 48.583 42.699 48.617 ;
      VIA 42.654 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 48.043 42.699 48.077 ;
      VIA 42.654 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 47.503 42.699 47.537 ;
      VIA 42.654 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 46.963 42.699 46.997 ;
      VIA 42.654 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 46.423 42.699 46.457 ;
      VIA 42.654 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 45.883 42.699 45.917 ;
      VIA 42.654 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 45.343 42.699 45.377 ;
      VIA 42.654 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 44.803 42.699 44.837 ;
      VIA 42.654 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 44.263 42.699 44.297 ;
      VIA 42.654 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 43.723 42.699 43.757 ;
      VIA 42.654 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 43.183 42.699 43.217 ;
      VIA 42.654 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 42.643 42.699 42.677 ;
      VIA 42.654 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 42.103 42.699 42.137 ;
      VIA 42.654 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 41.563 42.699 41.597 ;
      VIA 42.654 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 41.023 42.699 41.057 ;
      VIA 42.654 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 40.483 42.699 40.517 ;
      VIA 42.654 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 39.943 42.699 39.977 ;
      VIA 42.654 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 39.403 42.699 39.437 ;
      VIA 42.654 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 38.863 42.699 38.897 ;
      VIA 42.654 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 38.323 42.699 38.357 ;
      VIA 42.654 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 37.783 42.699 37.817 ;
      VIA 42.654 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 37.243 42.699 37.277 ;
      VIA 42.654 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 36.703 42.699 36.737 ;
      VIA 42.654 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 36.163 42.699 36.197 ;
      VIA 42.654 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 35.623 42.699 35.657 ;
      VIA 42.654 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 35.083 42.699 35.117 ;
      VIA 42.654 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 34.543 42.699 34.577 ;
      VIA 42.654 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 34.003 42.699 34.037 ;
      VIA 42.654 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 33.463 42.699 33.497 ;
      VIA 42.654 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 32.923 42.699 32.957 ;
      VIA 42.654 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 32.383 42.699 32.417 ;
      VIA 42.654 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 31.843 42.699 31.877 ;
      VIA 42.654 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 31.303 42.699 31.337 ;
      VIA 42.654 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 30.763 42.699 30.797 ;
      VIA 42.654 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 30.223 42.699 30.257 ;
      VIA 42.654 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 29.683 42.699 29.717 ;
      VIA 42.654 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 29.143 42.699 29.177 ;
      VIA 42.654 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 28.603 42.699 28.637 ;
      VIA 42.654 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 28.063 42.699 28.097 ;
      VIA 42.654 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 27.523 42.699 27.557 ;
      VIA 42.654 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 26.983 42.699 27.017 ;
      VIA 42.654 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 26.443 42.699 26.477 ;
      VIA 42.654 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 25.903 42.699 25.937 ;
      VIA 42.654 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 25.363 42.699 25.397 ;
      VIA 42.654 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 24.823 42.699 24.857 ;
      VIA 42.654 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 24.283 42.699 24.317 ;
      VIA 42.654 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 23.743 42.699 23.777 ;
      VIA 42.654 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 23.203 42.699 23.237 ;
      VIA 42.654 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 22.663 42.699 22.697 ;
      VIA 42.654 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 22.123 42.699 22.157 ;
      VIA 42.654 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 21.583 42.699 21.617 ;
      VIA 42.654 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 21.043 42.699 21.077 ;
      VIA 42.654 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 20.503 42.699 20.537 ;
      VIA 42.654 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 19.963 42.699 19.997 ;
      VIA 42.654 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 19.423 42.699 19.457 ;
      VIA 42.654 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 18.883 42.699 18.917 ;
      VIA 42.654 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 18.343 42.699 18.377 ;
      VIA 42.654 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 17.803 42.699 17.837 ;
      VIA 42.654 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 17.263 42.699 17.297 ;
      VIA 42.654 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 16.723 42.699 16.757 ;
      VIA 42.654 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 16.183 42.699 16.217 ;
      VIA 42.654 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 15.643 42.699 15.677 ;
      VIA 42.654 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 15.103 42.699 15.137 ;
      VIA 42.654 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 14.563 42.699 14.597 ;
      VIA 42.654 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 14.023 42.699 14.057 ;
      VIA 42.654 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 13.483 42.699 13.517 ;
      VIA 42.654 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 12.943 42.699 12.977 ;
      VIA 42.654 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 12.403 42.699 12.437 ;
      VIA 42.654 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 11.863 42.699 11.897 ;
      VIA 42.654 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 11.323 42.699 11.357 ;
      VIA 42.654 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 10.783 42.699 10.817 ;
      VIA 42.654 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 10.243 42.699 10.277 ;
      VIA 42.654 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 9.703 42.699 9.737 ;
      VIA 42.654 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 9.163 42.699 9.197 ;
      VIA 42.654 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 8.623 42.699 8.657 ;
      VIA 42.654 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 8.083 42.699 8.117 ;
      VIA 42.654 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 7.543 42.699 7.577 ;
      VIA 42.654 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 7.003 42.699 7.037 ;
      VIA 42.654 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 6.463 42.699 6.497 ;
      VIA 42.654 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 5.923 42.699 5.957 ;
      VIA 42.654 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 5.383 42.699 5.417 ;
      VIA 42.654 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 4.843 42.699 4.877 ;
      VIA 42.654 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 4.303 42.699 4.337 ;
      VIA 42.654 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 3.763 42.699 3.797 ;
      VIA 42.654 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 3.223 42.699 3.257 ;
      VIA 42.654 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 2.683 42.699 2.717 ;
      VIA 42.654 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 2.143 42.699 2.177 ;
      VIA 42.654 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 1.603 42.699 1.637 ;
      VIA 42.654 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 1.063 42.699 1.097 ;
      VIA 42.654 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 73.423 36.795 73.457 ;
      VIA 36.75 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 72.883 36.795 72.917 ;
      VIA 36.75 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 72.343 36.795 72.377 ;
      VIA 36.75 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 71.803 36.795 71.837 ;
      VIA 36.75 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 71.263 36.795 71.297 ;
      VIA 36.75 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 70.723 36.795 70.757 ;
      VIA 36.75 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 70.183 36.795 70.217 ;
      VIA 36.75 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 69.643 36.795 69.677 ;
      VIA 36.75 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 69.103 36.795 69.137 ;
      VIA 36.75 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 68.563 36.795 68.597 ;
      VIA 36.75 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 68.023 36.795 68.057 ;
      VIA 36.75 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 67.483 36.795 67.517 ;
      VIA 36.75 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 66.943 36.795 66.977 ;
      VIA 36.75 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 66.403 36.795 66.437 ;
      VIA 36.75 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 65.863 36.795 65.897 ;
      VIA 36.75 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 65.323 36.795 65.357 ;
      VIA 36.75 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 64.783 36.795 64.817 ;
      VIA 36.75 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 64.243 36.795 64.277 ;
      VIA 36.75 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 63.703 36.795 63.737 ;
      VIA 36.75 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 63.163 36.795 63.197 ;
      VIA 36.75 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 62.623 36.795 62.657 ;
      VIA 36.75 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 62.083 36.795 62.117 ;
      VIA 36.75 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 61.543 36.795 61.577 ;
      VIA 36.75 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 61.003 36.795 61.037 ;
      VIA 36.75 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 60.463 36.795 60.497 ;
      VIA 36.75 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 59.923 36.795 59.957 ;
      VIA 36.75 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 59.383 36.795 59.417 ;
      VIA 36.75 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 58.843 36.795 58.877 ;
      VIA 36.75 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 58.303 36.795 58.337 ;
      VIA 36.75 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 57.763 36.795 57.797 ;
      VIA 36.75 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 57.223 36.795 57.257 ;
      VIA 36.75 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 56.683 36.795 56.717 ;
      VIA 36.75 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 56.143 36.795 56.177 ;
      VIA 36.75 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 55.603 36.795 55.637 ;
      VIA 36.75 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 55.063 36.795 55.097 ;
      VIA 36.75 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 54.523 36.795 54.557 ;
      VIA 36.75 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 53.983 36.795 54.017 ;
      VIA 36.75 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 53.443 36.795 53.477 ;
      VIA 36.75 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 52.903 36.795 52.937 ;
      VIA 36.75 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 52.363 36.795 52.397 ;
      VIA 36.75 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 51.823 36.795 51.857 ;
      VIA 36.75 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 51.283 36.795 51.317 ;
      VIA 36.75 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 50.743 36.795 50.777 ;
      VIA 36.75 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 50.203 36.795 50.237 ;
      VIA 36.75 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 49.663 36.795 49.697 ;
      VIA 36.75 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 49.123 36.795 49.157 ;
      VIA 36.75 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 48.583 36.795 48.617 ;
      VIA 36.75 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 48.043 36.795 48.077 ;
      VIA 36.75 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 47.503 36.795 47.537 ;
      VIA 36.75 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 46.963 36.795 46.997 ;
      VIA 36.75 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 46.423 36.795 46.457 ;
      VIA 36.75 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 45.883 36.795 45.917 ;
      VIA 36.75 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 45.343 36.795 45.377 ;
      VIA 36.75 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 44.803 36.795 44.837 ;
      VIA 36.75 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 44.263 36.795 44.297 ;
      VIA 36.75 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 43.723 36.795 43.757 ;
      VIA 36.75 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 43.183 36.795 43.217 ;
      VIA 36.75 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 42.643 36.795 42.677 ;
      VIA 36.75 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 42.103 36.795 42.137 ;
      VIA 36.75 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 41.563 36.795 41.597 ;
      VIA 36.75 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 41.023 36.795 41.057 ;
      VIA 36.75 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 40.483 36.795 40.517 ;
      VIA 36.75 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.943 36.795 39.977 ;
      VIA 36.75 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.403 36.795 39.437 ;
      VIA 36.75 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.863 36.795 38.897 ;
      VIA 36.75 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.323 36.795 38.357 ;
      VIA 36.75 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.783 36.795 37.817 ;
      VIA 36.75 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.243 36.795 37.277 ;
      VIA 36.75 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.703 36.795 36.737 ;
      VIA 36.75 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.163 36.795 36.197 ;
      VIA 36.75 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.623 36.795 35.657 ;
      VIA 36.75 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.083 36.795 35.117 ;
      VIA 36.75 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.543 36.795 34.577 ;
      VIA 36.75 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.003 36.795 34.037 ;
      VIA 36.75 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 33.463 36.795 33.497 ;
      VIA 36.75 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.923 36.795 32.957 ;
      VIA 36.75 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.383 36.795 32.417 ;
      VIA 36.75 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.843 36.795 31.877 ;
      VIA 36.75 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.303 36.795 31.337 ;
      VIA 36.75 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.763 36.795 30.797 ;
      VIA 36.75 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.223 36.795 30.257 ;
      VIA 36.75 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.683 36.795 29.717 ;
      VIA 36.75 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.143 36.795 29.177 ;
      VIA 36.75 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.603 36.795 28.637 ;
      VIA 36.75 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.063 36.795 28.097 ;
      VIA 36.75 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 27.523 36.795 27.557 ;
      VIA 36.75 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.983 36.795 27.017 ;
      VIA 36.75 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.443 36.795 26.477 ;
      VIA 36.75 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.903 36.795 25.937 ;
      VIA 36.75 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.363 36.795 25.397 ;
      VIA 36.75 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.823 36.795 24.857 ;
      VIA 36.75 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.283 36.795 24.317 ;
      VIA 36.75 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.743 36.795 23.777 ;
      VIA 36.75 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.203 36.795 23.237 ;
      VIA 36.75 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.663 36.795 22.697 ;
      VIA 36.75 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.123 36.795 22.157 ;
      VIA 36.75 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.583 36.795 21.617 ;
      VIA 36.75 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.043 36.795 21.077 ;
      VIA 36.75 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 20.503 36.795 20.537 ;
      VIA 36.75 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.963 36.795 19.997 ;
      VIA 36.75 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.423 36.795 19.457 ;
      VIA 36.75 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.883 36.795 18.917 ;
      VIA 36.75 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.343 36.795 18.377 ;
      VIA 36.75 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.803 36.795 17.837 ;
      VIA 36.75 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.263 36.795 17.297 ;
      VIA 36.75 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.723 36.795 16.757 ;
      VIA 36.75 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.183 36.795 16.217 ;
      VIA 36.75 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.643 36.795 15.677 ;
      VIA 36.75 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.103 36.795 15.137 ;
      VIA 36.75 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.563 36.795 14.597 ;
      VIA 36.75 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.023 36.795 14.057 ;
      VIA 36.75 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 13.483 36.795 13.517 ;
      VIA 36.75 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.943 36.795 12.977 ;
      VIA 36.75 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.403 36.795 12.437 ;
      VIA 36.75 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.863 36.795 11.897 ;
      VIA 36.75 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.323 36.795 11.357 ;
      VIA 36.75 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.783 36.795 10.817 ;
      VIA 36.75 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.243 36.795 10.277 ;
      VIA 36.75 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.703 36.795 9.737 ;
      VIA 36.75 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.163 36.795 9.197 ;
      VIA 36.75 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.623 36.795 8.657 ;
      VIA 36.75 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.083 36.795 8.117 ;
      VIA 36.75 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.543 36.795 7.577 ;
      VIA 36.75 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.003 36.795 7.037 ;
      VIA 36.75 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 6.463 36.795 6.497 ;
      VIA 36.75 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.923 36.795 5.957 ;
      VIA 36.75 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.383 36.795 5.417 ;
      VIA 36.75 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.843 36.795 4.877 ;
      VIA 36.75 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.303 36.795 4.337 ;
      VIA 36.75 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.763 36.795 3.797 ;
      VIA 36.75 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.223 36.795 3.257 ;
      VIA 36.75 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.683 36.795 2.717 ;
      VIA 36.75 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.143 36.795 2.177 ;
      VIA 36.75 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.603 36.795 1.637 ;
      VIA 36.75 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.063 36.795 1.097 ;
      VIA 36.75 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 73.423 30.891 73.457 ;
      VIA 30.846 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 72.883 30.891 72.917 ;
      VIA 30.846 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 72.343 30.891 72.377 ;
      VIA 30.846 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 71.803 30.891 71.837 ;
      VIA 30.846 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 71.263 30.891 71.297 ;
      VIA 30.846 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 70.723 30.891 70.757 ;
      VIA 30.846 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 70.183 30.891 70.217 ;
      VIA 30.846 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 69.643 30.891 69.677 ;
      VIA 30.846 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 69.103 30.891 69.137 ;
      VIA 30.846 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 68.563 30.891 68.597 ;
      VIA 30.846 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 68.023 30.891 68.057 ;
      VIA 30.846 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 67.483 30.891 67.517 ;
      VIA 30.846 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 66.943 30.891 66.977 ;
      VIA 30.846 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 66.403 30.891 66.437 ;
      VIA 30.846 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 65.863 30.891 65.897 ;
      VIA 30.846 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 65.323 30.891 65.357 ;
      VIA 30.846 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 64.783 30.891 64.817 ;
      VIA 30.846 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 64.243 30.891 64.277 ;
      VIA 30.846 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 63.703 30.891 63.737 ;
      VIA 30.846 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 63.163 30.891 63.197 ;
      VIA 30.846 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 62.623 30.891 62.657 ;
      VIA 30.846 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 62.083 30.891 62.117 ;
      VIA 30.846 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 61.543 30.891 61.577 ;
      VIA 30.846 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 61.003 30.891 61.037 ;
      VIA 30.846 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 60.463 30.891 60.497 ;
      VIA 30.846 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 59.923 30.891 59.957 ;
      VIA 30.846 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 59.383 30.891 59.417 ;
      VIA 30.846 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 58.843 30.891 58.877 ;
      VIA 30.846 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 58.303 30.891 58.337 ;
      VIA 30.846 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 57.763 30.891 57.797 ;
      VIA 30.846 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 57.223 30.891 57.257 ;
      VIA 30.846 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 56.683 30.891 56.717 ;
      VIA 30.846 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 56.143 30.891 56.177 ;
      VIA 30.846 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 55.603 30.891 55.637 ;
      VIA 30.846 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 55.063 30.891 55.097 ;
      VIA 30.846 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 54.523 30.891 54.557 ;
      VIA 30.846 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 53.983 30.891 54.017 ;
      VIA 30.846 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 53.443 30.891 53.477 ;
      VIA 30.846 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 52.903 30.891 52.937 ;
      VIA 30.846 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 52.363 30.891 52.397 ;
      VIA 30.846 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 51.823 30.891 51.857 ;
      VIA 30.846 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 51.283 30.891 51.317 ;
      VIA 30.846 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 50.743 30.891 50.777 ;
      VIA 30.846 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 50.203 30.891 50.237 ;
      VIA 30.846 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 49.663 30.891 49.697 ;
      VIA 30.846 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 49.123 30.891 49.157 ;
      VIA 30.846 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 48.583 30.891 48.617 ;
      VIA 30.846 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 48.043 30.891 48.077 ;
      VIA 30.846 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 47.503 30.891 47.537 ;
      VIA 30.846 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 46.963 30.891 46.997 ;
      VIA 30.846 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 46.423 30.891 46.457 ;
      VIA 30.846 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 45.883 30.891 45.917 ;
      VIA 30.846 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 45.343 30.891 45.377 ;
      VIA 30.846 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 44.803 30.891 44.837 ;
      VIA 30.846 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 44.263 30.891 44.297 ;
      VIA 30.846 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 43.723 30.891 43.757 ;
      VIA 30.846 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 43.183 30.891 43.217 ;
      VIA 30.846 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 42.643 30.891 42.677 ;
      VIA 30.846 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 42.103 30.891 42.137 ;
      VIA 30.846 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 41.563 30.891 41.597 ;
      VIA 30.846 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 41.023 30.891 41.057 ;
      VIA 30.846 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 40.483 30.891 40.517 ;
      VIA 30.846 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.943 30.891 39.977 ;
      VIA 30.846 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.403 30.891 39.437 ;
      VIA 30.846 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.863 30.891 38.897 ;
      VIA 30.846 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.323 30.891 38.357 ;
      VIA 30.846 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.783 30.891 37.817 ;
      VIA 30.846 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.243 30.891 37.277 ;
      VIA 30.846 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.703 30.891 36.737 ;
      VIA 30.846 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.163 30.891 36.197 ;
      VIA 30.846 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.623 30.891 35.657 ;
      VIA 30.846 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.083 30.891 35.117 ;
      VIA 30.846 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.543 30.891 34.577 ;
      VIA 30.846 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.003 30.891 34.037 ;
      VIA 30.846 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 33.463 30.891 33.497 ;
      VIA 30.846 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.923 30.891 32.957 ;
      VIA 30.846 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.383 30.891 32.417 ;
      VIA 30.846 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.843 30.891 31.877 ;
      VIA 30.846 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.303 30.891 31.337 ;
      VIA 30.846 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.763 30.891 30.797 ;
      VIA 30.846 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.223 30.891 30.257 ;
      VIA 30.846 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.683 30.891 29.717 ;
      VIA 30.846 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.143 30.891 29.177 ;
      VIA 30.846 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.603 30.891 28.637 ;
      VIA 30.846 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.063 30.891 28.097 ;
      VIA 30.846 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 27.523 30.891 27.557 ;
      VIA 30.846 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.983 30.891 27.017 ;
      VIA 30.846 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.443 30.891 26.477 ;
      VIA 30.846 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.903 30.891 25.937 ;
      VIA 30.846 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.363 30.891 25.397 ;
      VIA 30.846 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.823 30.891 24.857 ;
      VIA 30.846 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.283 30.891 24.317 ;
      VIA 30.846 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.743 30.891 23.777 ;
      VIA 30.846 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.203 30.891 23.237 ;
      VIA 30.846 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.663 30.891 22.697 ;
      VIA 30.846 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.123 30.891 22.157 ;
      VIA 30.846 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.583 30.891 21.617 ;
      VIA 30.846 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.043 30.891 21.077 ;
      VIA 30.846 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 20.503 30.891 20.537 ;
      VIA 30.846 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.963 30.891 19.997 ;
      VIA 30.846 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.423 30.891 19.457 ;
      VIA 30.846 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.883 30.891 18.917 ;
      VIA 30.846 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.343 30.891 18.377 ;
      VIA 30.846 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.803 30.891 17.837 ;
      VIA 30.846 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.263 30.891 17.297 ;
      VIA 30.846 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.723 30.891 16.757 ;
      VIA 30.846 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.183 30.891 16.217 ;
      VIA 30.846 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.643 30.891 15.677 ;
      VIA 30.846 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.103 30.891 15.137 ;
      VIA 30.846 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.563 30.891 14.597 ;
      VIA 30.846 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.023 30.891 14.057 ;
      VIA 30.846 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 13.483 30.891 13.517 ;
      VIA 30.846 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.943 30.891 12.977 ;
      VIA 30.846 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.403 30.891 12.437 ;
      VIA 30.846 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.863 30.891 11.897 ;
      VIA 30.846 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.323 30.891 11.357 ;
      VIA 30.846 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.783 30.891 10.817 ;
      VIA 30.846 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.243 30.891 10.277 ;
      VIA 30.846 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.703 30.891 9.737 ;
      VIA 30.846 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.163 30.891 9.197 ;
      VIA 30.846 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.623 30.891 8.657 ;
      VIA 30.846 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.083 30.891 8.117 ;
      VIA 30.846 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.543 30.891 7.577 ;
      VIA 30.846 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.003 30.891 7.037 ;
      VIA 30.846 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 6.463 30.891 6.497 ;
      VIA 30.846 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.923 30.891 5.957 ;
      VIA 30.846 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.383 30.891 5.417 ;
      VIA 30.846 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.843 30.891 4.877 ;
      VIA 30.846 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.303 30.891 4.337 ;
      VIA 30.846 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.763 30.891 3.797 ;
      VIA 30.846 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.223 30.891 3.257 ;
      VIA 30.846 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.683 30.891 2.717 ;
      VIA 30.846 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.143 30.891 2.177 ;
      VIA 30.846 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.603 30.891 1.637 ;
      VIA 30.846 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.063 30.891 1.097 ;
      VIA 30.846 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 73.423 24.987 73.457 ;
      VIA 24.942 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 72.883 24.987 72.917 ;
      VIA 24.942 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 72.343 24.987 72.377 ;
      VIA 24.942 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 71.803 24.987 71.837 ;
      VIA 24.942 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 71.263 24.987 71.297 ;
      VIA 24.942 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 70.723 24.987 70.757 ;
      VIA 24.942 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 70.183 24.987 70.217 ;
      VIA 24.942 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 69.643 24.987 69.677 ;
      VIA 24.942 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 69.103 24.987 69.137 ;
      VIA 24.942 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 68.563 24.987 68.597 ;
      VIA 24.942 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 68.023 24.987 68.057 ;
      VIA 24.942 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 67.483 24.987 67.517 ;
      VIA 24.942 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 66.943 24.987 66.977 ;
      VIA 24.942 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 66.403 24.987 66.437 ;
      VIA 24.942 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 65.863 24.987 65.897 ;
      VIA 24.942 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 65.323 24.987 65.357 ;
      VIA 24.942 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 64.783 24.987 64.817 ;
      VIA 24.942 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 64.243 24.987 64.277 ;
      VIA 24.942 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 63.703 24.987 63.737 ;
      VIA 24.942 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 63.163 24.987 63.197 ;
      VIA 24.942 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 62.623 24.987 62.657 ;
      VIA 24.942 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 62.083 24.987 62.117 ;
      VIA 24.942 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 61.543 24.987 61.577 ;
      VIA 24.942 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 61.003 24.987 61.037 ;
      VIA 24.942 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 60.463 24.987 60.497 ;
      VIA 24.942 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 59.923 24.987 59.957 ;
      VIA 24.942 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 59.383 24.987 59.417 ;
      VIA 24.942 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 58.843 24.987 58.877 ;
      VIA 24.942 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 58.303 24.987 58.337 ;
      VIA 24.942 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 57.763 24.987 57.797 ;
      VIA 24.942 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 57.223 24.987 57.257 ;
      VIA 24.942 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 56.683 24.987 56.717 ;
      VIA 24.942 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 56.143 24.987 56.177 ;
      VIA 24.942 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 55.603 24.987 55.637 ;
      VIA 24.942 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 55.063 24.987 55.097 ;
      VIA 24.942 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 54.523 24.987 54.557 ;
      VIA 24.942 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 53.983 24.987 54.017 ;
      VIA 24.942 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 53.443 24.987 53.477 ;
      VIA 24.942 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 52.903 24.987 52.937 ;
      VIA 24.942 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 52.363 24.987 52.397 ;
      VIA 24.942 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 51.823 24.987 51.857 ;
      VIA 24.942 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 51.283 24.987 51.317 ;
      VIA 24.942 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 50.743 24.987 50.777 ;
      VIA 24.942 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 50.203 24.987 50.237 ;
      VIA 24.942 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 49.663 24.987 49.697 ;
      VIA 24.942 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 49.123 24.987 49.157 ;
      VIA 24.942 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 48.583 24.987 48.617 ;
      VIA 24.942 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 48.043 24.987 48.077 ;
      VIA 24.942 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 47.503 24.987 47.537 ;
      VIA 24.942 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 46.963 24.987 46.997 ;
      VIA 24.942 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 46.423 24.987 46.457 ;
      VIA 24.942 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 45.883 24.987 45.917 ;
      VIA 24.942 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 45.343 24.987 45.377 ;
      VIA 24.942 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 44.803 24.987 44.837 ;
      VIA 24.942 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 44.263 24.987 44.297 ;
      VIA 24.942 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 43.723 24.987 43.757 ;
      VIA 24.942 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 43.183 24.987 43.217 ;
      VIA 24.942 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 42.643 24.987 42.677 ;
      VIA 24.942 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 42.103 24.987 42.137 ;
      VIA 24.942 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 41.563 24.987 41.597 ;
      VIA 24.942 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 41.023 24.987 41.057 ;
      VIA 24.942 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 40.483 24.987 40.517 ;
      VIA 24.942 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.943 24.987 39.977 ;
      VIA 24.942 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.403 24.987 39.437 ;
      VIA 24.942 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.863 24.987 38.897 ;
      VIA 24.942 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.323 24.987 38.357 ;
      VIA 24.942 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.783 24.987 37.817 ;
      VIA 24.942 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.243 24.987 37.277 ;
      VIA 24.942 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.703 24.987 36.737 ;
      VIA 24.942 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.163 24.987 36.197 ;
      VIA 24.942 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.623 24.987 35.657 ;
      VIA 24.942 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.083 24.987 35.117 ;
      VIA 24.942 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.543 24.987 34.577 ;
      VIA 24.942 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.003 24.987 34.037 ;
      VIA 24.942 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 33.463 24.987 33.497 ;
      VIA 24.942 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.923 24.987 32.957 ;
      VIA 24.942 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.383 24.987 32.417 ;
      VIA 24.942 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.843 24.987 31.877 ;
      VIA 24.942 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.303 24.987 31.337 ;
      VIA 24.942 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.763 24.987 30.797 ;
      VIA 24.942 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.223 24.987 30.257 ;
      VIA 24.942 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.683 24.987 29.717 ;
      VIA 24.942 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.143 24.987 29.177 ;
      VIA 24.942 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.603 24.987 28.637 ;
      VIA 24.942 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.063 24.987 28.097 ;
      VIA 24.942 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 27.523 24.987 27.557 ;
      VIA 24.942 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.983 24.987 27.017 ;
      VIA 24.942 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.443 24.987 26.477 ;
      VIA 24.942 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.903 24.987 25.937 ;
      VIA 24.942 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.363 24.987 25.397 ;
      VIA 24.942 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.823 24.987 24.857 ;
      VIA 24.942 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.283 24.987 24.317 ;
      VIA 24.942 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.743 24.987 23.777 ;
      VIA 24.942 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.203 24.987 23.237 ;
      VIA 24.942 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.663 24.987 22.697 ;
      VIA 24.942 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.123 24.987 22.157 ;
      VIA 24.942 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.583 24.987 21.617 ;
      VIA 24.942 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.043 24.987 21.077 ;
      VIA 24.942 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 20.503 24.987 20.537 ;
      VIA 24.942 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.963 24.987 19.997 ;
      VIA 24.942 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.423 24.987 19.457 ;
      VIA 24.942 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.883 24.987 18.917 ;
      VIA 24.942 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.343 24.987 18.377 ;
      VIA 24.942 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.803 24.987 17.837 ;
      VIA 24.942 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.263 24.987 17.297 ;
      VIA 24.942 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.723 24.987 16.757 ;
      VIA 24.942 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.183 24.987 16.217 ;
      VIA 24.942 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.643 24.987 15.677 ;
      VIA 24.942 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.103 24.987 15.137 ;
      VIA 24.942 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.563 24.987 14.597 ;
      VIA 24.942 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.023 24.987 14.057 ;
      VIA 24.942 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 13.483 24.987 13.517 ;
      VIA 24.942 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.943 24.987 12.977 ;
      VIA 24.942 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.403 24.987 12.437 ;
      VIA 24.942 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.863 24.987 11.897 ;
      VIA 24.942 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.323 24.987 11.357 ;
      VIA 24.942 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.783 24.987 10.817 ;
      VIA 24.942 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.243 24.987 10.277 ;
      VIA 24.942 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.703 24.987 9.737 ;
      VIA 24.942 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.163 24.987 9.197 ;
      VIA 24.942 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.623 24.987 8.657 ;
      VIA 24.942 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.083 24.987 8.117 ;
      VIA 24.942 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.543 24.987 7.577 ;
      VIA 24.942 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.003 24.987 7.037 ;
      VIA 24.942 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 6.463 24.987 6.497 ;
      VIA 24.942 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.923 24.987 5.957 ;
      VIA 24.942 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.383 24.987 5.417 ;
      VIA 24.942 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.843 24.987 4.877 ;
      VIA 24.942 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.303 24.987 4.337 ;
      VIA 24.942 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.763 24.987 3.797 ;
      VIA 24.942 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.223 24.987 3.257 ;
      VIA 24.942 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.683 24.987 2.717 ;
      VIA 24.942 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.143 24.987 2.177 ;
      VIA 24.942 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.603 24.987 1.637 ;
      VIA 24.942 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.063 24.987 1.097 ;
      VIA 24.942 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 73.423 19.083 73.457 ;
      VIA 19.038 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 72.883 19.083 72.917 ;
      VIA 19.038 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 72.343 19.083 72.377 ;
      VIA 19.038 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 71.803 19.083 71.837 ;
      VIA 19.038 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 71.263 19.083 71.297 ;
      VIA 19.038 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 70.723 19.083 70.757 ;
      VIA 19.038 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 70.183 19.083 70.217 ;
      VIA 19.038 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 69.643 19.083 69.677 ;
      VIA 19.038 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 69.103 19.083 69.137 ;
      VIA 19.038 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 68.563 19.083 68.597 ;
      VIA 19.038 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 68.023 19.083 68.057 ;
      VIA 19.038 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 67.483 19.083 67.517 ;
      VIA 19.038 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 66.943 19.083 66.977 ;
      VIA 19.038 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 66.403 19.083 66.437 ;
      VIA 19.038 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 65.863 19.083 65.897 ;
      VIA 19.038 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 65.323 19.083 65.357 ;
      VIA 19.038 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 64.783 19.083 64.817 ;
      VIA 19.038 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 64.243 19.083 64.277 ;
      VIA 19.038 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 63.703 19.083 63.737 ;
      VIA 19.038 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 63.163 19.083 63.197 ;
      VIA 19.038 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 62.623 19.083 62.657 ;
      VIA 19.038 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 62.083 19.083 62.117 ;
      VIA 19.038 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 61.543 19.083 61.577 ;
      VIA 19.038 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 61.003 19.083 61.037 ;
      VIA 19.038 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 60.463 19.083 60.497 ;
      VIA 19.038 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 59.923 19.083 59.957 ;
      VIA 19.038 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 59.383 19.083 59.417 ;
      VIA 19.038 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 58.843 19.083 58.877 ;
      VIA 19.038 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 58.303 19.083 58.337 ;
      VIA 19.038 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 57.763 19.083 57.797 ;
      VIA 19.038 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 57.223 19.083 57.257 ;
      VIA 19.038 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 56.683 19.083 56.717 ;
      VIA 19.038 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 56.143 19.083 56.177 ;
      VIA 19.038 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 55.603 19.083 55.637 ;
      VIA 19.038 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 55.063 19.083 55.097 ;
      VIA 19.038 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 54.523 19.083 54.557 ;
      VIA 19.038 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 53.983 19.083 54.017 ;
      VIA 19.038 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 53.443 19.083 53.477 ;
      VIA 19.038 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 52.903 19.083 52.937 ;
      VIA 19.038 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 52.363 19.083 52.397 ;
      VIA 19.038 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 51.823 19.083 51.857 ;
      VIA 19.038 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 51.283 19.083 51.317 ;
      VIA 19.038 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 50.743 19.083 50.777 ;
      VIA 19.038 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 50.203 19.083 50.237 ;
      VIA 19.038 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 49.663 19.083 49.697 ;
      VIA 19.038 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 49.123 19.083 49.157 ;
      VIA 19.038 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 48.583 19.083 48.617 ;
      VIA 19.038 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 48.043 19.083 48.077 ;
      VIA 19.038 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 47.503 19.083 47.537 ;
      VIA 19.038 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 46.963 19.083 46.997 ;
      VIA 19.038 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 46.423 19.083 46.457 ;
      VIA 19.038 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 45.883 19.083 45.917 ;
      VIA 19.038 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 45.343 19.083 45.377 ;
      VIA 19.038 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 44.803 19.083 44.837 ;
      VIA 19.038 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 44.263 19.083 44.297 ;
      VIA 19.038 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 43.723 19.083 43.757 ;
      VIA 19.038 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 43.183 19.083 43.217 ;
      VIA 19.038 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 42.643 19.083 42.677 ;
      VIA 19.038 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 42.103 19.083 42.137 ;
      VIA 19.038 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 41.563 19.083 41.597 ;
      VIA 19.038 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 41.023 19.083 41.057 ;
      VIA 19.038 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 40.483 19.083 40.517 ;
      VIA 19.038 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.943 19.083 39.977 ;
      VIA 19.038 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.403 19.083 39.437 ;
      VIA 19.038 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.863 19.083 38.897 ;
      VIA 19.038 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.323 19.083 38.357 ;
      VIA 19.038 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.783 19.083 37.817 ;
      VIA 19.038 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.243 19.083 37.277 ;
      VIA 19.038 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.703 19.083 36.737 ;
      VIA 19.038 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.163 19.083 36.197 ;
      VIA 19.038 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.623 19.083 35.657 ;
      VIA 19.038 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.083 19.083 35.117 ;
      VIA 19.038 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.543 19.083 34.577 ;
      VIA 19.038 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.003 19.083 34.037 ;
      VIA 19.038 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 33.463 19.083 33.497 ;
      VIA 19.038 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.923 19.083 32.957 ;
      VIA 19.038 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.383 19.083 32.417 ;
      VIA 19.038 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.843 19.083 31.877 ;
      VIA 19.038 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.303 19.083 31.337 ;
      VIA 19.038 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.763 19.083 30.797 ;
      VIA 19.038 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.223 19.083 30.257 ;
      VIA 19.038 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.683 19.083 29.717 ;
      VIA 19.038 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.143 19.083 29.177 ;
      VIA 19.038 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.603 19.083 28.637 ;
      VIA 19.038 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.063 19.083 28.097 ;
      VIA 19.038 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 27.523 19.083 27.557 ;
      VIA 19.038 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.983 19.083 27.017 ;
      VIA 19.038 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.443 19.083 26.477 ;
      VIA 19.038 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.903 19.083 25.937 ;
      VIA 19.038 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.363 19.083 25.397 ;
      VIA 19.038 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.823 19.083 24.857 ;
      VIA 19.038 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.283 19.083 24.317 ;
      VIA 19.038 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.743 19.083 23.777 ;
      VIA 19.038 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.203 19.083 23.237 ;
      VIA 19.038 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.663 19.083 22.697 ;
      VIA 19.038 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.123 19.083 22.157 ;
      VIA 19.038 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.583 19.083 21.617 ;
      VIA 19.038 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.043 19.083 21.077 ;
      VIA 19.038 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 20.503 19.083 20.537 ;
      VIA 19.038 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.963 19.083 19.997 ;
      VIA 19.038 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.423 19.083 19.457 ;
      VIA 19.038 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.883 19.083 18.917 ;
      VIA 19.038 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.343 19.083 18.377 ;
      VIA 19.038 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.803 19.083 17.837 ;
      VIA 19.038 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.263 19.083 17.297 ;
      VIA 19.038 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.723 19.083 16.757 ;
      VIA 19.038 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.183 19.083 16.217 ;
      VIA 19.038 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.643 19.083 15.677 ;
      VIA 19.038 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.103 19.083 15.137 ;
      VIA 19.038 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.563 19.083 14.597 ;
      VIA 19.038 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.023 19.083 14.057 ;
      VIA 19.038 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 13.483 19.083 13.517 ;
      VIA 19.038 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.943 19.083 12.977 ;
      VIA 19.038 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.403 19.083 12.437 ;
      VIA 19.038 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.863 19.083 11.897 ;
      VIA 19.038 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.323 19.083 11.357 ;
      VIA 19.038 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.783 19.083 10.817 ;
      VIA 19.038 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.243 19.083 10.277 ;
      VIA 19.038 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.703 19.083 9.737 ;
      VIA 19.038 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.163 19.083 9.197 ;
      VIA 19.038 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.623 19.083 8.657 ;
      VIA 19.038 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.083 19.083 8.117 ;
      VIA 19.038 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.543 19.083 7.577 ;
      VIA 19.038 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.003 19.083 7.037 ;
      VIA 19.038 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 6.463 19.083 6.497 ;
      VIA 19.038 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.923 19.083 5.957 ;
      VIA 19.038 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.383 19.083 5.417 ;
      VIA 19.038 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.843 19.083 4.877 ;
      VIA 19.038 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.303 19.083 4.337 ;
      VIA 19.038 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.763 19.083 3.797 ;
      VIA 19.038 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.223 19.083 3.257 ;
      VIA 19.038 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.683 19.083 2.717 ;
      VIA 19.038 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.143 19.083 2.177 ;
      VIA 19.038 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.603 19.083 1.637 ;
      VIA 19.038 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.063 19.083 1.097 ;
      VIA 19.038 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 73.423 13.179 73.457 ;
      VIA 13.134 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 72.883 13.179 72.917 ;
      VIA 13.134 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 72.343 13.179 72.377 ;
      VIA 13.134 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 71.803 13.179 71.837 ;
      VIA 13.134 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 71.263 13.179 71.297 ;
      VIA 13.134 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 70.723 13.179 70.757 ;
      VIA 13.134 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 70.183 13.179 70.217 ;
      VIA 13.134 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 69.643 13.179 69.677 ;
      VIA 13.134 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 69.103 13.179 69.137 ;
      VIA 13.134 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 68.563 13.179 68.597 ;
      VIA 13.134 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 68.023 13.179 68.057 ;
      VIA 13.134 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 67.483 13.179 67.517 ;
      VIA 13.134 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 66.943 13.179 66.977 ;
      VIA 13.134 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 66.403 13.179 66.437 ;
      VIA 13.134 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 65.863 13.179 65.897 ;
      VIA 13.134 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 65.323 13.179 65.357 ;
      VIA 13.134 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 64.783 13.179 64.817 ;
      VIA 13.134 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 64.243 13.179 64.277 ;
      VIA 13.134 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 63.703 13.179 63.737 ;
      VIA 13.134 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 63.163 13.179 63.197 ;
      VIA 13.134 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 62.623 13.179 62.657 ;
      VIA 13.134 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 62.083 13.179 62.117 ;
      VIA 13.134 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 61.543 13.179 61.577 ;
      VIA 13.134 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 61.003 13.179 61.037 ;
      VIA 13.134 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 60.463 13.179 60.497 ;
      VIA 13.134 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 59.923 13.179 59.957 ;
      VIA 13.134 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 59.383 13.179 59.417 ;
      VIA 13.134 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 58.843 13.179 58.877 ;
      VIA 13.134 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 58.303 13.179 58.337 ;
      VIA 13.134 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 57.763 13.179 57.797 ;
      VIA 13.134 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 57.223 13.179 57.257 ;
      VIA 13.134 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 56.683 13.179 56.717 ;
      VIA 13.134 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 56.143 13.179 56.177 ;
      VIA 13.134 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 55.603 13.179 55.637 ;
      VIA 13.134 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 55.063 13.179 55.097 ;
      VIA 13.134 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 54.523 13.179 54.557 ;
      VIA 13.134 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 53.983 13.179 54.017 ;
      VIA 13.134 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 53.443 13.179 53.477 ;
      VIA 13.134 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 52.903 13.179 52.937 ;
      VIA 13.134 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 52.363 13.179 52.397 ;
      VIA 13.134 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 51.823 13.179 51.857 ;
      VIA 13.134 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 51.283 13.179 51.317 ;
      VIA 13.134 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 50.743 13.179 50.777 ;
      VIA 13.134 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 50.203 13.179 50.237 ;
      VIA 13.134 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 49.663 13.179 49.697 ;
      VIA 13.134 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 49.123 13.179 49.157 ;
      VIA 13.134 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 48.583 13.179 48.617 ;
      VIA 13.134 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 48.043 13.179 48.077 ;
      VIA 13.134 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 47.503 13.179 47.537 ;
      VIA 13.134 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 46.963 13.179 46.997 ;
      VIA 13.134 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 46.423 13.179 46.457 ;
      VIA 13.134 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 45.883 13.179 45.917 ;
      VIA 13.134 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 45.343 13.179 45.377 ;
      VIA 13.134 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 44.803 13.179 44.837 ;
      VIA 13.134 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 44.263 13.179 44.297 ;
      VIA 13.134 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 43.723 13.179 43.757 ;
      VIA 13.134 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 43.183 13.179 43.217 ;
      VIA 13.134 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 42.643 13.179 42.677 ;
      VIA 13.134 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 42.103 13.179 42.137 ;
      VIA 13.134 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 41.563 13.179 41.597 ;
      VIA 13.134 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 41.023 13.179 41.057 ;
      VIA 13.134 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 40.483 13.179 40.517 ;
      VIA 13.134 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.943 13.179 39.977 ;
      VIA 13.134 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.403 13.179 39.437 ;
      VIA 13.134 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.863 13.179 38.897 ;
      VIA 13.134 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.323 13.179 38.357 ;
      VIA 13.134 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.783 13.179 37.817 ;
      VIA 13.134 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.243 13.179 37.277 ;
      VIA 13.134 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.703 13.179 36.737 ;
      VIA 13.134 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.163 13.179 36.197 ;
      VIA 13.134 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.623 13.179 35.657 ;
      VIA 13.134 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.083 13.179 35.117 ;
      VIA 13.134 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.543 13.179 34.577 ;
      VIA 13.134 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.003 13.179 34.037 ;
      VIA 13.134 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 33.463 13.179 33.497 ;
      VIA 13.134 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.923 13.179 32.957 ;
      VIA 13.134 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.383 13.179 32.417 ;
      VIA 13.134 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.843 13.179 31.877 ;
      VIA 13.134 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.303 13.179 31.337 ;
      VIA 13.134 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.763 13.179 30.797 ;
      VIA 13.134 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.223 13.179 30.257 ;
      VIA 13.134 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.683 13.179 29.717 ;
      VIA 13.134 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.143 13.179 29.177 ;
      VIA 13.134 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.603 13.179 28.637 ;
      VIA 13.134 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.063 13.179 28.097 ;
      VIA 13.134 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 27.523 13.179 27.557 ;
      VIA 13.134 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.983 13.179 27.017 ;
      VIA 13.134 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.443 13.179 26.477 ;
      VIA 13.134 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.903 13.179 25.937 ;
      VIA 13.134 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.363 13.179 25.397 ;
      VIA 13.134 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.823 13.179 24.857 ;
      VIA 13.134 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.283 13.179 24.317 ;
      VIA 13.134 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.743 13.179 23.777 ;
      VIA 13.134 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.203 13.179 23.237 ;
      VIA 13.134 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.663 13.179 22.697 ;
      VIA 13.134 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.123 13.179 22.157 ;
      VIA 13.134 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.583 13.179 21.617 ;
      VIA 13.134 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.043 13.179 21.077 ;
      VIA 13.134 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 20.503 13.179 20.537 ;
      VIA 13.134 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.963 13.179 19.997 ;
      VIA 13.134 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.423 13.179 19.457 ;
      VIA 13.134 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.883 13.179 18.917 ;
      VIA 13.134 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.343 13.179 18.377 ;
      VIA 13.134 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.803 13.179 17.837 ;
      VIA 13.134 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.263 13.179 17.297 ;
      VIA 13.134 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.723 13.179 16.757 ;
      VIA 13.134 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.183 13.179 16.217 ;
      VIA 13.134 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.643 13.179 15.677 ;
      VIA 13.134 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.103 13.179 15.137 ;
      VIA 13.134 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.563 13.179 14.597 ;
      VIA 13.134 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.023 13.179 14.057 ;
      VIA 13.134 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 13.483 13.179 13.517 ;
      VIA 13.134 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.943 13.179 12.977 ;
      VIA 13.134 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.403 13.179 12.437 ;
      VIA 13.134 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.863 13.179 11.897 ;
      VIA 13.134 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.323 13.179 11.357 ;
      VIA 13.134 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.783 13.179 10.817 ;
      VIA 13.134 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.243 13.179 10.277 ;
      VIA 13.134 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.703 13.179 9.737 ;
      VIA 13.134 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.163 13.179 9.197 ;
      VIA 13.134 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.623 13.179 8.657 ;
      VIA 13.134 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.083 13.179 8.117 ;
      VIA 13.134 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.543 13.179 7.577 ;
      VIA 13.134 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.003 13.179 7.037 ;
      VIA 13.134 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 6.463 13.179 6.497 ;
      VIA 13.134 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.923 13.179 5.957 ;
      VIA 13.134 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.383 13.179 5.417 ;
      VIA 13.134 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.843 13.179 4.877 ;
      VIA 13.134 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.303 13.179 4.337 ;
      VIA 13.134 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.763 13.179 3.797 ;
      VIA 13.134 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.223 13.179 3.257 ;
      VIA 13.134 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.683 13.179 2.717 ;
      VIA 13.134 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.143 13.179 2.177 ;
      VIA 13.134 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.603 13.179 1.637 ;
      VIA 13.134 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.063 13.179 1.097 ;
      VIA 13.134 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 73.423 7.275 73.457 ;
      VIA 7.23 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 72.883 7.275 72.917 ;
      VIA 7.23 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 72.343 7.275 72.377 ;
      VIA 7.23 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 71.803 7.275 71.837 ;
      VIA 7.23 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 71.263 7.275 71.297 ;
      VIA 7.23 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 70.723 7.275 70.757 ;
      VIA 7.23 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 70.183 7.275 70.217 ;
      VIA 7.23 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 69.643 7.275 69.677 ;
      VIA 7.23 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 69.103 7.275 69.137 ;
      VIA 7.23 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 68.563 7.275 68.597 ;
      VIA 7.23 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 68.023 7.275 68.057 ;
      VIA 7.23 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 67.483 7.275 67.517 ;
      VIA 7.23 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 66.943 7.275 66.977 ;
      VIA 7.23 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 66.403 7.275 66.437 ;
      VIA 7.23 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 65.863 7.275 65.897 ;
      VIA 7.23 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 65.323 7.275 65.357 ;
      VIA 7.23 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 64.783 7.275 64.817 ;
      VIA 7.23 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 64.243 7.275 64.277 ;
      VIA 7.23 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 63.703 7.275 63.737 ;
      VIA 7.23 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 63.163 7.275 63.197 ;
      VIA 7.23 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 62.623 7.275 62.657 ;
      VIA 7.23 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 62.083 7.275 62.117 ;
      VIA 7.23 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 61.543 7.275 61.577 ;
      VIA 7.23 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 61.003 7.275 61.037 ;
      VIA 7.23 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 60.463 7.275 60.497 ;
      VIA 7.23 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 59.923 7.275 59.957 ;
      VIA 7.23 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 59.383 7.275 59.417 ;
      VIA 7.23 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 58.843 7.275 58.877 ;
      VIA 7.23 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 58.303 7.275 58.337 ;
      VIA 7.23 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 57.763 7.275 57.797 ;
      VIA 7.23 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 57.223 7.275 57.257 ;
      VIA 7.23 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 56.683 7.275 56.717 ;
      VIA 7.23 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 56.143 7.275 56.177 ;
      VIA 7.23 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 55.603 7.275 55.637 ;
      VIA 7.23 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 55.063 7.275 55.097 ;
      VIA 7.23 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 54.523 7.275 54.557 ;
      VIA 7.23 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 53.983 7.275 54.017 ;
      VIA 7.23 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 53.443 7.275 53.477 ;
      VIA 7.23 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 52.903 7.275 52.937 ;
      VIA 7.23 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 52.363 7.275 52.397 ;
      VIA 7.23 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 51.823 7.275 51.857 ;
      VIA 7.23 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 51.283 7.275 51.317 ;
      VIA 7.23 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 50.743 7.275 50.777 ;
      VIA 7.23 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 50.203 7.275 50.237 ;
      VIA 7.23 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 49.663 7.275 49.697 ;
      VIA 7.23 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 49.123 7.275 49.157 ;
      VIA 7.23 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 48.583 7.275 48.617 ;
      VIA 7.23 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 48.043 7.275 48.077 ;
      VIA 7.23 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 47.503 7.275 47.537 ;
      VIA 7.23 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 46.963 7.275 46.997 ;
      VIA 7.23 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 46.423 7.275 46.457 ;
      VIA 7.23 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 45.883 7.275 45.917 ;
      VIA 7.23 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 45.343 7.275 45.377 ;
      VIA 7.23 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 44.803 7.275 44.837 ;
      VIA 7.23 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 44.263 7.275 44.297 ;
      VIA 7.23 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 43.723 7.275 43.757 ;
      VIA 7.23 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 43.183 7.275 43.217 ;
      VIA 7.23 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 42.643 7.275 42.677 ;
      VIA 7.23 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 42.103 7.275 42.137 ;
      VIA 7.23 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 41.563 7.275 41.597 ;
      VIA 7.23 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 41.023 7.275 41.057 ;
      VIA 7.23 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 40.483 7.275 40.517 ;
      VIA 7.23 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.943 7.275 39.977 ;
      VIA 7.23 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.403 7.275 39.437 ;
      VIA 7.23 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.863 7.275 38.897 ;
      VIA 7.23 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.323 7.275 38.357 ;
      VIA 7.23 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.783 7.275 37.817 ;
      VIA 7.23 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.243 7.275 37.277 ;
      VIA 7.23 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.703 7.275 36.737 ;
      VIA 7.23 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.163 7.275 36.197 ;
      VIA 7.23 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.623 7.275 35.657 ;
      VIA 7.23 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.083 7.275 35.117 ;
      VIA 7.23 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.543 7.275 34.577 ;
      VIA 7.23 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.003 7.275 34.037 ;
      VIA 7.23 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 33.463 7.275 33.497 ;
      VIA 7.23 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.923 7.275 32.957 ;
      VIA 7.23 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.383 7.275 32.417 ;
      VIA 7.23 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.843 7.275 31.877 ;
      VIA 7.23 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.303 7.275 31.337 ;
      VIA 7.23 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.763 7.275 30.797 ;
      VIA 7.23 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.223 7.275 30.257 ;
      VIA 7.23 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.683 7.275 29.717 ;
      VIA 7.23 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.143 7.275 29.177 ;
      VIA 7.23 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.603 7.275 28.637 ;
      VIA 7.23 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.063 7.275 28.097 ;
      VIA 7.23 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 27.523 7.275 27.557 ;
      VIA 7.23 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.983 7.275 27.017 ;
      VIA 7.23 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.443 7.275 26.477 ;
      VIA 7.23 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.903 7.275 25.937 ;
      VIA 7.23 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.363 7.275 25.397 ;
      VIA 7.23 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.823 7.275 24.857 ;
      VIA 7.23 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.283 7.275 24.317 ;
      VIA 7.23 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.743 7.275 23.777 ;
      VIA 7.23 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.203 7.275 23.237 ;
      VIA 7.23 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.663 7.275 22.697 ;
      VIA 7.23 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.123 7.275 22.157 ;
      VIA 7.23 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.583 7.275 21.617 ;
      VIA 7.23 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.043 7.275 21.077 ;
      VIA 7.23 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 20.503 7.275 20.537 ;
      VIA 7.23 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.963 7.275 19.997 ;
      VIA 7.23 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.423 7.275 19.457 ;
      VIA 7.23 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.883 7.275 18.917 ;
      VIA 7.23 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.343 7.275 18.377 ;
      VIA 7.23 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.803 7.275 17.837 ;
      VIA 7.23 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.263 7.275 17.297 ;
      VIA 7.23 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.723 7.275 16.757 ;
      VIA 7.23 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.183 7.275 16.217 ;
      VIA 7.23 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.643 7.275 15.677 ;
      VIA 7.23 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.103 7.275 15.137 ;
      VIA 7.23 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.563 7.275 14.597 ;
      VIA 7.23 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.023 7.275 14.057 ;
      VIA 7.23 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 13.483 7.275 13.517 ;
      VIA 7.23 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.943 7.275 12.977 ;
      VIA 7.23 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.403 7.275 12.437 ;
      VIA 7.23 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.863 7.275 11.897 ;
      VIA 7.23 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.323 7.275 11.357 ;
      VIA 7.23 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.783 7.275 10.817 ;
      VIA 7.23 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.243 7.275 10.277 ;
      VIA 7.23 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.703 7.275 9.737 ;
      VIA 7.23 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.163 7.275 9.197 ;
      VIA 7.23 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.623 7.275 8.657 ;
      VIA 7.23 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.083 7.275 8.117 ;
      VIA 7.23 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.543 7.275 7.577 ;
      VIA 7.23 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.003 7.275 7.037 ;
      VIA 7.23 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 6.463 7.275 6.497 ;
      VIA 7.23 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.923 7.275 5.957 ;
      VIA 7.23 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.383 7.275 5.417 ;
      VIA 7.23 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.843 7.275 4.877 ;
      VIA 7.23 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.303 7.275 4.337 ;
      VIA 7.23 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.763 7.275 3.797 ;
      VIA 7.23 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.223 7.275 3.257 ;
      VIA 7.23 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.683 7.275 2.717 ;
      VIA 7.23 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.143 7.275 2.177 ;
      VIA 7.23 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.603 7.275 1.637 ;
      VIA 7.23 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.063 7.275 1.097 ;
      VIA 7.23 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 73.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 73.423 1.371 73.457 ;
      VIA 1.326 73.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 73.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 72.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 72.883 1.371 72.917 ;
      VIA 1.326 72.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 72.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 72.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 72.343 1.371 72.377 ;
      VIA 1.326 72.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 72.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 71.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 71.803 1.371 71.837 ;
      VIA 1.326 71.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 71.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 71.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 71.263 1.371 71.297 ;
      VIA 1.326 71.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 71.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 70.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 70.723 1.371 70.757 ;
      VIA 1.326 70.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 70.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 70.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 70.183 1.371 70.217 ;
      VIA 1.326 70.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 70.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 69.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 69.643 1.371 69.677 ;
      VIA 1.326 69.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 69.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 69.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 69.103 1.371 69.137 ;
      VIA 1.326 69.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 69.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 68.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 68.563 1.371 68.597 ;
      VIA 1.326 68.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 68.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 68.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 68.023 1.371 68.057 ;
      VIA 1.326 68.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 68.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 67.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 67.483 1.371 67.517 ;
      VIA 1.326 67.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 67.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 66.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 66.943 1.371 66.977 ;
      VIA 1.326 66.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 66.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 66.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 66.403 1.371 66.437 ;
      VIA 1.326 66.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 66.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 65.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 65.863 1.371 65.897 ;
      VIA 1.326 65.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 65.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 65.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 65.323 1.371 65.357 ;
      VIA 1.326 65.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 65.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 64.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 64.783 1.371 64.817 ;
      VIA 1.326 64.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 64.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 64.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 64.243 1.371 64.277 ;
      VIA 1.326 64.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 64.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 63.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 63.703 1.371 63.737 ;
      VIA 1.326 63.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 63.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 63.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 63.163 1.371 63.197 ;
      VIA 1.326 63.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 63.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 62.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 62.623 1.371 62.657 ;
      VIA 1.326 62.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 62.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 62.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 62.083 1.371 62.117 ;
      VIA 1.326 62.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 62.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 61.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 61.543 1.371 61.577 ;
      VIA 1.326 61.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 61.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 61.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 61.003 1.371 61.037 ;
      VIA 1.326 61.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 61.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 60.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 60.463 1.371 60.497 ;
      VIA 1.326 60.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 60.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 59.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 59.923 1.371 59.957 ;
      VIA 1.326 59.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 59.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 59.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 59.383 1.371 59.417 ;
      VIA 1.326 59.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 59.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 58.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 58.843 1.371 58.877 ;
      VIA 1.326 58.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 58.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 58.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 58.303 1.371 58.337 ;
      VIA 1.326 58.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 58.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 57.763 1.371 57.797 ;
      VIA 1.326 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 57.223 1.371 57.257 ;
      VIA 1.326 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 56.683 1.371 56.717 ;
      VIA 1.326 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 56.143 1.371 56.177 ;
      VIA 1.326 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 55.603 1.371 55.637 ;
      VIA 1.326 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 55.063 1.371 55.097 ;
      VIA 1.326 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 54.523 1.371 54.557 ;
      VIA 1.326 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 53.983 1.371 54.017 ;
      VIA 1.326 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 53.443 1.371 53.477 ;
      VIA 1.326 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 52.903 1.371 52.937 ;
      VIA 1.326 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 52.363 1.371 52.397 ;
      VIA 1.326 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 51.823 1.371 51.857 ;
      VIA 1.326 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 51.283 1.371 51.317 ;
      VIA 1.326 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 50.743 1.371 50.777 ;
      VIA 1.326 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 50.203 1.371 50.237 ;
      VIA 1.326 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 49.663 1.371 49.697 ;
      VIA 1.326 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 49.123 1.371 49.157 ;
      VIA 1.326 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 48.583 1.371 48.617 ;
      VIA 1.326 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 48.043 1.371 48.077 ;
      VIA 1.326 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 47.503 1.371 47.537 ;
      VIA 1.326 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 46.963 1.371 46.997 ;
      VIA 1.326 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 46.423 1.371 46.457 ;
      VIA 1.326 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 45.883 1.371 45.917 ;
      VIA 1.326 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 45.343 1.371 45.377 ;
      VIA 1.326 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 44.803 1.371 44.837 ;
      VIA 1.326 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 44.263 1.371 44.297 ;
      VIA 1.326 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 43.723 1.371 43.757 ;
      VIA 1.326 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 43.183 1.371 43.217 ;
      VIA 1.326 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 42.643 1.371 42.677 ;
      VIA 1.326 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 42.103 1.371 42.137 ;
      VIA 1.326 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 41.563 1.371 41.597 ;
      VIA 1.326 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 41.023 1.371 41.057 ;
      VIA 1.326 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 40.483 1.371 40.517 ;
      VIA 1.326 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.943 1.371 39.977 ;
      VIA 1.326 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.403 1.371 39.437 ;
      VIA 1.326 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.863 1.371 38.897 ;
      VIA 1.326 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.323 1.371 38.357 ;
      VIA 1.326 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.783 1.371 37.817 ;
      VIA 1.326 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.243 1.371 37.277 ;
      VIA 1.326 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.703 1.371 36.737 ;
      VIA 1.326 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.163 1.371 36.197 ;
      VIA 1.326 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.623 1.371 35.657 ;
      VIA 1.326 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.083 1.371 35.117 ;
      VIA 1.326 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.543 1.371 34.577 ;
      VIA 1.326 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.003 1.371 34.037 ;
      VIA 1.326 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 33.463 1.371 33.497 ;
      VIA 1.326 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.923 1.371 32.957 ;
      VIA 1.326 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.383 1.371 32.417 ;
      VIA 1.326 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.843 1.371 31.877 ;
      VIA 1.326 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.303 1.371 31.337 ;
      VIA 1.326 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.763 1.371 30.797 ;
      VIA 1.326 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.223 1.371 30.257 ;
      VIA 1.326 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.683 1.371 29.717 ;
      VIA 1.326 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.143 1.371 29.177 ;
      VIA 1.326 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.603 1.371 28.637 ;
      VIA 1.326 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.063 1.371 28.097 ;
      VIA 1.326 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 27.523 1.371 27.557 ;
      VIA 1.326 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.983 1.371 27.017 ;
      VIA 1.326 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.443 1.371 26.477 ;
      VIA 1.326 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.903 1.371 25.937 ;
      VIA 1.326 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.363 1.371 25.397 ;
      VIA 1.326 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.823 1.371 24.857 ;
      VIA 1.326 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.283 1.371 24.317 ;
      VIA 1.326 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.743 1.371 23.777 ;
      VIA 1.326 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.203 1.371 23.237 ;
      VIA 1.326 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.663 1.371 22.697 ;
      VIA 1.326 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.123 1.371 22.157 ;
      VIA 1.326 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.583 1.371 21.617 ;
      VIA 1.326 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.043 1.371 21.077 ;
      VIA 1.326 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 20.503 1.371 20.537 ;
      VIA 1.326 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.963 1.371 19.997 ;
      VIA 1.326 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.423 1.371 19.457 ;
      VIA 1.326 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.883 1.371 18.917 ;
      VIA 1.326 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.343 1.371 18.377 ;
      VIA 1.326 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.803 1.371 17.837 ;
      VIA 1.326 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.263 1.371 17.297 ;
      VIA 1.326 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.723 1.371 16.757 ;
      VIA 1.326 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.183 1.371 16.217 ;
      VIA 1.326 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.643 1.371 15.677 ;
      VIA 1.326 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.103 1.371 15.137 ;
      VIA 1.326 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.563 1.371 14.597 ;
      VIA 1.326 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.023 1.371 14.057 ;
      VIA 1.326 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 13.483 1.371 13.517 ;
      VIA 1.326 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.943 1.371 12.977 ;
      VIA 1.326 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.403 1.371 12.437 ;
      VIA 1.326 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.863 1.371 11.897 ;
      VIA 1.326 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.323 1.371 11.357 ;
      VIA 1.326 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.783 1.371 10.817 ;
      VIA 1.326 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.243 1.371 10.277 ;
      VIA 1.326 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.703 1.371 9.737 ;
      VIA 1.326 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.163 1.371 9.197 ;
      VIA 1.326 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.623 1.371 8.657 ;
      VIA 1.326 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.083 1.371 8.117 ;
      VIA 1.326 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.543 1.371 7.577 ;
      VIA 1.326 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.003 1.371 7.037 ;
      VIA 1.326 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 6.463 1.371 6.497 ;
      VIA 1.326 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.923 1.371 5.957 ;
      VIA 1.326 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.383 1.371 5.417 ;
      VIA 1.326 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 37.341 73.44 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 72.9 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 72.36 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 71.82 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 71.28 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 70.74 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 70.2 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 69.66 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 69.12 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 68.58 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 68.04 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 67.5 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 66.96 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 66.42 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 65.88 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 65.34 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 64.8 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 64.26 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 63.72 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 63.18 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 62.64 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 62.1 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 61.56 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 61.02 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 60.48 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 59.94 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 59.4 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 58.86 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 58.32 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 57.78 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 57.24 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 56.7 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 56.16 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 55.62 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 55.08 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 54.54 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 54 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 53.46 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 52.92 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 52.38 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 51.84 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 51.3 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 50.76 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 50.22 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 49.68 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 49.14 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 48.6 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 48.06 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 47.52 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 46.98 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 46.44 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 45.9 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 45.36 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 44.82 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 44.28 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 43.74 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 43.2 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 42.66 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 42.12 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 41.58 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 41.04 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 40.5 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 39.96 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 39.42 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 38.88 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 38.34 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 37.8 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 37.26 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 36.72 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 36.18 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 35.64 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 35.1 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 34.56 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 34.02 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 33.48 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 32.94 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 32.4 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 31.86 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 31.32 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 30.78 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 30.24 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 29.7 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 29.16 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 28.62 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 28.08 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 27.54 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 27 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 26.46 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 25.92 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 25.38 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 24.84 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 24.3 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 23.76 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 23.22 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 22.68 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 22.14 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 21.6 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 21.06 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 20.52 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 19.98 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 19.44 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 18.9 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 18.36 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 17.82 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 17.28 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 16.74 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 16.2 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 15.66 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 15.12 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 14.58 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 14.04 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 13.5 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 12.96 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 12.42 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 11.88 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 11.34 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 10.8 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 10.26 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 9.72 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 9.18 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 8.64 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 8.1 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 7.56 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 7.02 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 6.48 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 5.94 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 5.4 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 4.86 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 4.32 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 3.78 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 3.24 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 2.7 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 2.16 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 1.62 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
      VIA 37.341 1.08 run_benchmark_via1_2_72630_18_1_2017_36_36 ;
    END
  END VSS
  PIN M_DataRdy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.672 0 0.696 0.084 ;
    END
  END M_DataRdy[0]
  PIN M_DataRdy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.768 0 0.792 0.084 ;
    END
  END M_DataRdy[1]
  PIN M_Rdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 39.456 0.084 39.48 ;
    END
  END M_Rdata_ram[0]
  PIN M_Rdata_ram[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.752 74.707 34.776 ;
    END
  END M_Rdata_ram[100]
  PIN M_Rdata_ram[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.52 74.707 35.544 ;
    END
  END M_Rdata_ram[101]
  PIN M_Rdata_ram[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.36 74.707 39.384 ;
    END
  END M_Rdata_ram[102]
  PIN M_Rdata_ram[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.128 74.707 52.152 ;
    END
  END M_Rdata_ram[103]
  PIN M_Rdata_ram[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.264 74.707 39.288 ;
    END
  END M_Rdata_ram[104]
  PIN M_Rdata_ram[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.616 74.707 35.64 ;
    END
  END M_Rdata_ram[105]
  PIN M_Rdata_ram[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.136 74.707 35.16 ;
    END
  END M_Rdata_ram[106]
  PIN M_Rdata_ram[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.936 74.707 39.96 ;
    END
  END M_Rdata_ram[107]
  PIN M_Rdata_ram[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.84 74.707 39.864 ;
    END
  END M_Rdata_ram[108]
  PIN M_Rdata_ram[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.744 74.707 39.768 ;
    END
  END M_Rdata_ram[109]
  PIN M_Rdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 38.4 0.084 38.424 ;
    END
  END M_Rdata_ram[10]
  PIN M_Rdata_ram[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.4 74.707 38.424 ;
    END
  END M_Rdata_ram[110]
  PIN M_Rdata_ram[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.76 74.707 41.784 ;
    END
  END M_Rdata_ram[111]
  PIN M_Rdata_ram[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.552 74.707 39.576 ;
    END
  END M_Rdata_ram[112]
  PIN M_Rdata_ram[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.456 74.707 39.48 ;
    END
  END M_Rdata_ram[113]
  PIN M_Rdata_ram[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.512 74.707 40.536 ;
    END
  END M_Rdata_ram[114]
  PIN M_Rdata_ram[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.088 74.707 41.112 ;
    END
  END M_Rdata_ram[115]
  PIN M_Rdata_ram[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.08 74.707 46.104 ;
    END
  END M_Rdata_ram[116]
  PIN M_Rdata_ram[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.04 74.707 47.064 ;
    END
  END M_Rdata_ram[117]
  PIN M_Rdata_ram[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.008 74.707 43.032 ;
    END
  END M_Rdata_ram[118]
  PIN M_Rdata_ram[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.528 74.707 42.552 ;
    END
  END M_Rdata_ram[119]
  PIN M_Rdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 40.128 0.084 40.152 ;
    END
  END M_Rdata_ram[11]
  PIN M_Rdata_ram[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.52 74.707 47.544 ;
    END
  END M_Rdata_ram[120]
  PIN M_Rdata_ram[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.424 74.707 47.448 ;
    END
  END M_Rdata_ram[121]
  PIN M_Rdata_ram[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.328 74.707 47.352 ;
    END
  END M_Rdata_ram[122]
  PIN M_Rdata_ram[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.312 74.707 45.336 ;
    END
  END M_Rdata_ram[123]
  PIN M_Rdata_ram[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.736 74.707 44.76 ;
    END
  END M_Rdata_ram[124]
  PIN M_Rdata_ram[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.68 74.707 43.704 ;
    END
  END M_Rdata_ram[125]
  PIN M_Rdata_ram[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.584 74.707 43.608 ;
    END
  END M_Rdata_ram[126]
  PIN M_Rdata_ram[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.928 74.707 44.952 ;
    END
  END M_Rdata_ram[127]
  PIN M_Rdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 41.28 0.084 41.304 ;
    END
  END M_Rdata_ram[12]
  PIN M_Rdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 40.608 0.084 40.632 ;
    END
  END M_Rdata_ram[13]
  PIN M_Rdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 42.144 0.084 42.168 ;
    END
  END M_Rdata_ram[14]
  PIN M_Rdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 40.512 0.084 40.536 ;
    END
  END M_Rdata_ram[15]
  PIN M_Rdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 39.36 0.084 39.384 ;
    END
  END M_Rdata_ram[16]
  PIN M_Rdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 38.016 0.084 38.04 ;
    END
  END M_Rdata_ram[17]
  PIN M_Rdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 38.112 0.084 38.136 ;
    END
  END M_Rdata_ram[18]
  PIN M_Rdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 39.168 0.084 39.192 ;
    END
  END M_Rdata_ram[19]
  PIN M_Rdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 38.688 0.084 38.712 ;
    END
  END M_Rdata_ram[1]
  PIN M_Rdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 34.848 0.084 34.872 ;
    END
  END M_Rdata_ram[20]
  PIN M_Rdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 35.52 0.084 35.544 ;
    END
  END M_Rdata_ram[21]
  PIN M_Rdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 34.944 0.084 34.968 ;
    END
  END M_Rdata_ram[22]
  PIN M_Rdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 34.752 0.084 34.776 ;
    END
  END M_Rdata_ram[23]
  PIN M_Rdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.432 0.084 30.456 ;
    END
  END M_Rdata_ram[24]
  PIN M_Rdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.856 0.084 29.88 ;
    END
  END M_Rdata_ram[25]
  PIN M_Rdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.952 0.084 29.976 ;
    END
  END M_Rdata_ram[26]
  PIN M_Rdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.144 0.084 30.168 ;
    END
  END M_Rdata_ram[27]
  PIN M_Rdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.568 0.084 29.592 ;
    END
  END M_Rdata_ram[28]
  PIN M_Rdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.896 0.084 28.92 ;
    END
  END M_Rdata_ram[29]
  PIN M_Rdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 39.264 0.084 39.288 ;
    END
  END M_Rdata_ram[2]
  PIN M_Rdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.8 0.084 28.824 ;
    END
  END M_Rdata_ram[30]
  PIN M_Rdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.992 0.084 29.016 ;
    END
  END M_Rdata_ram[31]
  PIN M_Rdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 41.952 0.084 41.976 ;
    END
  END M_Rdata_ram[32]
  PIN M_Rdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 42.24 0.084 42.264 ;
    END
  END M_Rdata_ram[33]
  PIN M_Rdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 42.048 0.084 42.072 ;
    END
  END M_Rdata_ram[34]
  PIN M_Rdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 43.2 0.084 43.224 ;
    END
  END M_Rdata_ram[35]
  PIN M_Rdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 42.912 0.084 42.936 ;
    END
  END M_Rdata_ram[36]
  PIN M_Rdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 43.776 0.084 43.8 ;
    END
  END M_Rdata_ram[37]
  PIN M_Rdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 43.008 0.084 43.032 ;
    END
  END M_Rdata_ram[38]
  PIN M_Rdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 44.448 0.084 44.472 ;
    END
  END M_Rdata_ram[39]
  PIN M_Rdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 38.88 0.084 38.904 ;
    END
  END M_Rdata_ram[3]
  PIN M_Rdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.504 0.084 45.528 ;
    END
  END M_Rdata_ram[40]
  PIN M_Rdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 46.368 0.084 46.392 ;
    END
  END M_Rdata_ram[41]
  PIN M_Rdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.216 0.084 45.24 ;
    END
  END M_Rdata_ram[42]
  PIN M_Rdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.6 0.084 45.624 ;
    END
  END M_Rdata_ram[43]
  PIN M_Rdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 43.968 0.084 43.992 ;
    END
  END M_Rdata_ram[44]
  PIN M_Rdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 44.352 0.084 44.376 ;
    END
  END M_Rdata_ram[45]
  PIN M_Rdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 43.872 0.084 43.896 ;
    END
  END M_Rdata_ram[46]
  PIN M_Rdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 44.256 0.084 44.28 ;
    END
  END M_Rdata_ram[47]
  PIN M_Rdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.12 0.084 45.144 ;
    END
  END M_Rdata_ram[48]
  PIN M_Rdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.024 0.084 45.048 ;
    END
  END M_Rdata_ram[49]
  PIN M_Rdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.728 0.084 37.752 ;
    END
  END M_Rdata_ram[4]
  PIN M_Rdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 45.792 0.084 45.816 ;
    END
  END M_Rdata_ram[50]
  PIN M_Rdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 46.752 0.084 46.776 ;
    END
  END M_Rdata_ram[51]
  PIN M_Rdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.616 74.623 47.64 74.707 ;
    END
  END M_Rdata_ram[52]
  PIN M_Rdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.52 74.623 47.544 74.707 ;
    END
  END M_Rdata_ram[53]
  PIN M_Rdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.808 74.623 47.832 74.707 ;
    END
  END M_Rdata_ram[54]
  PIN M_Rdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.424 74.623 47.448 74.707 ;
    END
  END M_Rdata_ram[55]
  PIN M_Rdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.328 74.623 47.352 74.707 ;
    END
  END M_Rdata_ram[56]
  PIN M_Rdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  47.712 74.623 47.736 74.707 ;
    END
  END M_Rdata_ram[57]
  PIN M_Rdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  48 74.623 48.024 74.707 ;
    END
  END M_Rdata_ram[58]
  PIN M_Rdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  49.44 74.623 49.464 74.707 ;
    END
  END M_Rdata_ram[59]
  PIN M_Rdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.152 0.084 37.176 ;
    END
  END M_Rdata_ram[5]
  PIN M_Rdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  49.056 74.623 49.08 74.707 ;
    END
  END M_Rdata_ram[60]
  PIN M_Rdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  50.304 74.623 50.328 74.707 ;
    END
  END M_Rdata_ram[61]
  PIN M_Rdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  50.016 74.623 50.04 74.707 ;
    END
  END M_Rdata_ram[62]
  PIN M_Rdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.456 74.707 51.48 ;
    END
  END M_Rdata_ram[63]
  PIN M_Rdata_ram[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.752 74.707 46.776 ;
    END
  END M_Rdata_ram[64]
  PIN M_Rdata_ram[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.656 74.707 46.68 ;
    END
  END M_Rdata_ram[65]
  PIN M_Rdata_ram[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.504 74.707 45.528 ;
    END
  END M_Rdata_ram[66]
  PIN M_Rdata_ram[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.464 74.707 46.488 ;
    END
  END M_Rdata_ram[67]
  PIN M_Rdata_ram[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.368 74.707 46.392 ;
    END
  END M_Rdata_ram[68]
  PIN M_Rdata_ram[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.56 74.707 46.584 ;
    END
  END M_Rdata_ram[69]
  PIN M_Rdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.248 0.084 37.272 ;
    END
  END M_Rdata_ram[6]
  PIN M_Rdata_ram[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.272 74.707 46.296 ;
    END
  END M_Rdata_ram[70]
  PIN M_Rdata_ram[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.232 74.707 47.256 ;
    END
  END M_Rdata_ram[71]
  PIN M_Rdata_ram[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.136 74.707 47.16 ;
    END
  END M_Rdata_ram[72]
  PIN M_Rdata_ram[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.288 74.707 48.312 ;
    END
  END M_Rdata_ram[73]
  PIN M_Rdata_ram[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.264 74.707 51.288 ;
    END
  END M_Rdata_ram[74]
  PIN M_Rdata_ram[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.248 74.707 49.272 ;
    END
  END M_Rdata_ram[75]
  PIN M_Rdata_ram[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.688 74.707 50.712 ;
    END
  END M_Rdata_ram[76]
  PIN M_Rdata_ram[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.112 74.707 50.136 ;
    END
  END M_Rdata_ram[77]
  PIN M_Rdata_ram[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.4 74.707 50.424 ;
    END
  END M_Rdata_ram[78]
  PIN M_Rdata_ram[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.496 74.707 50.52 ;
    END
  END M_Rdata_ram[79]
  PIN M_Rdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.056 0.084 37.08 ;
    END
  END M_Rdata_ram[7]
  PIN M_Rdata_ram[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.536 74.707 49.56 ;
    END
  END M_Rdata_ram[80]
  PIN M_Rdata_ram[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.92 74.707 49.944 ;
    END
  END M_Rdata_ram[81]
  PIN M_Rdata_ram[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.304 74.707 50.328 ;
    END
  END M_Rdata_ram[82]
  PIN M_Rdata_ram[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.88 74.707 50.904 ;
    END
  END M_Rdata_ram[83]
  PIN M_Rdata_ram[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.544 74.707 32.568 ;
    END
  END M_Rdata_ram[84]
  PIN M_Rdata_ram[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 30.912 74.707 30.936 ;
    END
  END M_Rdata_ram[85]
  PIN M_Rdata_ram[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.392 74.707 31.416 ;
    END
  END M_Rdata_ram[86]
  PIN M_Rdata_ram[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.216 74.707 33.24 ;
    END
  END M_Rdata_ram[87]
  PIN M_Rdata_ram[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.504 74.707 33.528 ;
    END
  END M_Rdata_ram[88]
  PIN M_Rdata_ram[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.928 74.707 32.952 ;
    END
  END M_Rdata_ram[89]
  PIN M_Rdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 39.072 0.084 39.096 ;
    END
  END M_Rdata_ram[8]
  PIN M_Rdata_ram[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.984 74.707 34.008 ;
    END
  END M_Rdata_ram[90]
  PIN M_Rdata_ram[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.464 74.707 34.488 ;
    END
  END M_Rdata_ram[91]
  PIN M_Rdata_ram[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.096 74.707 36.12 ;
    END
  END M_Rdata_ram[92]
  PIN M_Rdata_ram[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36 74.707 36.024 ;
    END
  END M_Rdata_ram[93]
  PIN M_Rdata_ram[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.344 74.707 37.368 ;
    END
  END M_Rdata_ram[94]
  PIN M_Rdata_ram[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.384 74.707 36.408 ;
    END
  END M_Rdata_ram[95]
  PIN M_Rdata_ram[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.48 74.707 36.504 ;
    END
  END M_Rdata_ram[96]
  PIN M_Rdata_ram[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.424 74.707 35.448 ;
    END
  END M_Rdata_ram[97]
  PIN M_Rdata_ram[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.04 74.707 35.064 ;
    END
  END M_Rdata_ram[98]
  PIN M_Rdata_ram[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.728 74.707 37.752 ;
    END
  END M_Rdata_ram[99]
  PIN M_Rdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.92 0.084 37.944 ;
    END
  END M_Rdata_ram[9]
  PIN Min_Wdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.632 74.707 37.656 ;
    END
  END Min_Wdata_ram[0]
  PIN Min_Wdata_ram[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.376 74.623 53.4 74.707 ;
    END
  END Min_Wdata_ram[100]
  PIN Min_Wdata_ram[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.864 74.623 60.888 74.707 ;
    END
  END Min_Wdata_ram[101]
  PIN Min_Wdata_ram[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.648 0.084 3.672 ;
    END
  END Min_Wdata_ram[102]
  PIN Min_Wdata_ram[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.56 74.623 58.584 74.707 ;
    END
  END Min_Wdata_ram[103]
  PIN Min_Wdata_ram[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.536 74.623 13.56 74.707 ;
    END
  END Min_Wdata_ram[104]
  PIN Min_Wdata_ram[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.024 74.623 33.048 74.707 ;
    END
  END Min_Wdata_ram[105]
  PIN Min_Wdata_ram[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.368 0 58.392 0.084 ;
    END
  END Min_Wdata_ram[106]
  PIN Min_Wdata_ram[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.04 0 59.064 0.084 ;
    END
  END Min_Wdata_ram[107]
  PIN Min_Wdata_ram[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.624 74.623 6.648 74.707 ;
    END
  END Min_Wdata_ram[108]
  PIN Min_Wdata_ram[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.968 0 31.992 0.084 ;
    END
  END Min_Wdata_ram[109]
  PIN Min_Wdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.44 74.707 37.464 ;
    END
  END Min_Wdata_ram[10]
  PIN Min_Wdata_ram[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.856 0 53.88 0.084 ;
    END
  END Min_Wdata_ram[110]
  PIN Min_Wdata_ram[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.344 0 61.368 0.084 ;
    END
  END Min_Wdata_ram[111]
  PIN Min_Wdata_ram[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.4 0 62.424 0.084 ;
    END
  END Min_Wdata_ram[112]
  PIN Min_Wdata_ram[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 70.656 74.707 70.68 ;
    END
  END Min_Wdata_ram[113]
  PIN Min_Wdata_ram[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.176 74.623 34.2 74.707 ;
    END
  END Min_Wdata_ram[114]
  PIN Min_Wdata_ram[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.168 0 63.192 0.084 ;
    END
  END Min_Wdata_ram[115]
  PIN Min_Wdata_ram[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.328 74.623 59.352 74.707 ;
    END
  END Min_Wdata_ram[116]
  PIN Min_Wdata_ram[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.504 74.623 57.528 74.707 ;
    END
  END Min_Wdata_ram[117]
  PIN Min_Wdata_ram[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.92 74.623 37.944 74.707 ;
    END
  END Min_Wdata_ram[118]
  PIN Min_Wdata_ram[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.6 74.623 57.624 74.707 ;
    END
  END Min_Wdata_ram[119]
  PIN Min_Wdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.688 74.707 38.712 ;
    END
  END Min_Wdata_ram[11]
  PIN Min_Wdata_ram[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.688 0 62.712 0.084 ;
    END
  END Min_Wdata_ram[120]
  PIN Min_Wdata_ram[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.472 74.623 41.496 74.707 ;
    END
  END Min_Wdata_ram[121]
  PIN Min_Wdata_ram[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.168 0 39.192 0.084 ;
    END
  END Min_Wdata_ram[122]
  PIN Min_Wdata_ram[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.992 74.623 53.016 74.707 ;
    END
  END Min_Wdata_ram[123]
  PIN Min_Wdata_ram[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.44 0 61.464 0.084 ;
    END
  END Min_Wdata_ram[124]
  PIN Min_Wdata_ram[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.72 0 6.744 0.084 ;
    END
  END Min_Wdata_ram[125]
  PIN Min_Wdata_ram[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.576 0 36.6 0.084 ;
    END
  END Min_Wdata_ram[126]
  PIN Min_Wdata_ram[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.152 0 61.176 0.084 ;
    END
  END Min_Wdata_ram[127]
  PIN Min_Wdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.232 74.707 35.256 ;
    END
  END Min_Wdata_ram[12]
  PIN Min_Wdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.848 74.707 34.872 ;
    END
  END Min_Wdata_ram[13]
  PIN Min_Wdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.08 74.707 34.104 ;
    END
  END Min_Wdata_ram[14]
  PIN Min_Wdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.352 74.707 32.376 ;
    END
  END Min_Wdata_ram[15]
  PIN Min_Wdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.448 74.707 32.472 ;
    END
  END Min_Wdata_ram[16]
  PIN Min_Wdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.488 74.707 31.512 ;
    END
  END Min_Wdata_ram[17]
  PIN Min_Wdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.872 74.707 31.896 ;
    END
  END Min_Wdata_ram[18]
  PIN Min_Wdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.2 74.707 31.224 ;
    END
  END Min_Wdata_ram[19]
  PIN Min_Wdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.248 74.707 37.272 ;
    END
  END Min_Wdata_ram[1]
  PIN Min_Wdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.584 74.707 31.608 ;
    END
  END Min_Wdata_ram[20]
  PIN Min_Wdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.104 74.707 31.128 ;
    END
  END Min_Wdata_ram[21]
  PIN Min_Wdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.296 74.707 31.32 ;
    END
  END Min_Wdata_ram[22]
  PIN Min_Wdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.12 74.707 33.144 ;
    END
  END Min_Wdata_ram[23]
  PIN Min_Wdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.6 74.707 33.624 ;
    END
  END Min_Wdata_ram[24]
  PIN Min_Wdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.736 74.707 32.76 ;
    END
  END Min_Wdata_ram[25]
  PIN Min_Wdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.176 74.707 34.2 ;
    END
  END Min_Wdata_ram[26]
  PIN Min_Wdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.56 74.707 34.584 ;
    END
  END Min_Wdata_ram[27]
  PIN Min_Wdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.288 74.707 36.312 ;
    END
  END Min_Wdata_ram[28]
  PIN Min_Wdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.576 74.707 36.6 ;
    END
  END Min_Wdata_ram[29]
  PIN Min_Wdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.152 74.707 37.176 ;
    END
  END Min_Wdata_ram[2]
  PIN Min_Wdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.904 74.707 35.928 ;
    END
  END Min_Wdata_ram[30]
  PIN Min_Wdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.992 74.707 41.016 ;
    END
  END Min_Wdata_ram[31]
  PIN Min_Wdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.704 74.707 40.728 ;
    END
  END Min_Wdata_ram[32]
  PIN Min_Wdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  46.464 74.623 46.488 74.707 ;
    END
  END Min_Wdata_ram[33]
  PIN Min_Wdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.168 74.707 39.192 ;
    END
  END Min_Wdata_ram[34]
  PIN Min_Wdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.048 74.707 42.072 ;
    END
  END Min_Wdata_ram[35]
  PIN Min_Wdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.2 74.707 43.224 ;
    END
  END Min_Wdata_ram[36]
  PIN Min_Wdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.624 74.707 42.648 ;
    END
  END Min_Wdata_ram[37]
  PIN Min_Wdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.984 74.707 58.008 ;
    END
  END Min_Wdata_ram[38]
  PIN Min_Wdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.376 74.707 41.4 ;
    END
  END Min_Wdata_ram[39]
  PIN Min_Wdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.808 74.707 35.832 ;
    END
  END Min_Wdata_ram[3]
  PIN Min_Wdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.224 74.707 52.248 ;
    END
  END Min_Wdata_ram[40]
  PIN Min_Wdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.28 74.707 41.304 ;
    END
  END Min_Wdata_ram[41]
  PIN Min_Wdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.072 74.707 39.096 ;
    END
  END Min_Wdata_ram[42]
  PIN Min_Wdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.336 74.707 42.36 ;
    END
  END Min_Wdata_ram[43]
  PIN Min_Wdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.064 74.707 44.088 ;
    END
  END Min_Wdata_ram[44]
  PIN Min_Wdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.184 74.707 41.208 ;
    END
  END Min_Wdata_ram[45]
  PIN Min_Wdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.896 74.707 40.92 ;
    END
  END Min_Wdata_ram[46]
  PIN Min_Wdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.816 74.707 42.84 ;
    END
  END Min_Wdata_ram[47]
  PIN Min_Wdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.12 74.707 57.144 ;
    END
  END Min_Wdata_ram[48]
  PIN Min_Wdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.488 74.707 43.512 ;
    END
  END Min_Wdata_ram[49]
  PIN Min_Wdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.432 74.707 42.456 ;
    END
  END Min_Wdata_ram[4]
  PIN Min_Wdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.472 74.707 41.496 ;
    END
  END Min_Wdata_ram[50]
  PIN Min_Wdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.64 74.707 44.664 ;
    END
  END Min_Wdata_ram[51]
  PIN Min_Wdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.24 74.707 42.264 ;
    END
  END Min_Wdata_ram[52]
  PIN Min_Wdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.984 74.707 46.008 ;
    END
  END Min_Wdata_ram[53]
  PIN Min_Wdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.912 74.707 42.936 ;
    END
  END Min_Wdata_ram[54]
  PIN Min_Wdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.968 74.707 43.992 ;
    END
  END Min_Wdata_ram[55]
  PIN Min_Wdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.176 74.707 46.2 ;
    END
  END Min_Wdata_ram[56]
  PIN Min_Wdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.792 74.707 45.816 ;
    END
  END Min_Wdata_ram[57]
  PIN Min_Wdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.6 74.707 45.624 ;
    END
  END Min_Wdata_ram[58]
  PIN Min_Wdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.216 74.707 45.24 ;
    END
  END Min_Wdata_ram[59]
  PIN Min_Wdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.712 74.707 35.736 ;
    END
  END Min_Wdata_ram[5]
  PIN Min_Wdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.208 74.707 50.232 ;
    END
  END Min_Wdata_ram[60]
  PIN Min_Wdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.544 74.707 44.568 ;
    END
  END Min_Wdata_ram[61]
  PIN Min_Wdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.848 74.707 46.872 ;
    END
  END Min_Wdata_ram[62]
  PIN Min_Wdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.448 74.707 44.472 ;
    END
  END Min_Wdata_ram[63]
  PIN Min_Wdata_ram[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.944 74.623 22.968 74.707 ;
    END
  END Min_Wdata_ram[64]
  PIN Min_Wdata_ram[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.656 74.623 58.68 74.707 ;
    END
  END Min_Wdata_ram[65]
  PIN Min_Wdata_ram[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.752 74.623 58.776 74.707 ;
    END
  END Min_Wdata_ram[66]
  PIN Min_Wdata_ram[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  43.968 74.623 43.992 74.707 ;
    END
  END Min_Wdata_ram[67]
  PIN Min_Wdata_ram[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.56 0 34.584 0.084 ;
    END
  END Min_Wdata_ram[68]
  PIN Min_Wdata_ram[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.096 74.623 60.12 74.707 ;
    END
  END Min_Wdata_ram[69]
  PIN Min_Wdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.448 74.707 56.472 ;
    END
  END Min_Wdata_ram[6]
  PIN Min_Wdata_ram[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  66.624 74.623 66.648 74.707 ;
    END
  END Min_Wdata_ram[70]
  PIN Min_Wdata_ram[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  45.12 0 45.144 0.084 ;
    END
  END Min_Wdata_ram[71]
  PIN Min_Wdata_ram[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.288 74.623 60.312 74.707 ;
    END
  END Min_Wdata_ram[72]
  PIN Min_Wdata_ram[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.496 74.623 2.52 74.707 ;
    END
  END Min_Wdata_ram[73]
  PIN Min_Wdata_ram[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.28 74.623 53.304 74.707 ;
    END
  END Min_Wdata_ram[74]
  PIN Min_Wdata_ram[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.136 74.623 59.16 74.707 ;
    END
  END Min_Wdata_ram[75]
  PIN Min_Wdata_ram[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.184 0 17.208 0.084 ;
    END
  END Min_Wdata_ram[76]
  PIN Min_Wdata_ram[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.608 0 52.632 0.084 ;
    END
  END Min_Wdata_ram[77]
  PIN Min_Wdata_ram[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.608 74.623 52.632 74.707 ;
    END
  END Min_Wdata_ram[78]
  PIN Min_Wdata_ram[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.232 74.623 59.256 74.707 ;
    END
  END Min_Wdata_ram[79]
  PIN Min_Wdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.592 74.707 38.616 ;
    END
  END Min_Wdata_ram[7]
  PIN Min_Wdata_ram[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.624 74.623 54.648 74.707 ;
    END
  END Min_Wdata_ram[80]
  PIN Min_Wdata_ram[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.776 74.623 55.8 74.707 ;
    END
  END Min_Wdata_ram[81]
  PIN Min_Wdata_ram[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.464 0 34.488 0.084 ;
    END
  END Min_Wdata_ram[82]
  PIN Min_Wdata_ram[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.76 74.623 53.784 74.707 ;
    END
  END Min_Wdata_ram[83]
  PIN Min_Wdata_ram[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.384 0 60.408 0.084 ;
    END
  END Min_Wdata_ram[84]
  PIN Min_Wdata_ram[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.096 0 60.12 0.084 ;
    END
  END Min_Wdata_ram[85]
  PIN Min_Wdata_ram[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.216 74.623 21.24 74.707 ;
    END
  END Min_Wdata_ram[86]
  PIN Min_Wdata_ram[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  43.008 0 43.032 0.084 ;
    END
  END Min_Wdata_ram[87]
  PIN Min_Wdata_ram[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.04 74.623 59.064 74.707 ;
    END
  END Min_Wdata_ram[88]
  PIN Min_Wdata_ram[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 62.88 74.707 62.904 ;
    END
  END Min_Wdata_ram[89]
  PIN Min_Wdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.92 74.707 37.944 ;
    END
  END Min_Wdata_ram[8]
  PIN Min_Wdata_ram[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  45.504 74.623 45.528 74.707 ;
    END
  END Min_Wdata_ram[90]
  PIN Min_Wdata_ram[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.28 74.623 41.304 74.707 ;
    END
  END Min_Wdata_ram[91]
  PIN Min_Wdata_ram[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.072 0 39.096 0.084 ;
    END
  END Min_Wdata_ram[92]
  PIN Min_Wdata_ram[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.456 0 63.48 0.084 ;
    END
  END Min_Wdata_ram[93]
  PIN Min_Wdata_ram[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.416 74.623 52.44 74.707 ;
    END
  END Min_Wdata_ram[94]
  PIN Min_Wdata_ram[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.888 74.623 57.912 74.707 ;
    END
  END Min_Wdata_ram[95]
  PIN Min_Wdata_ram[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.48 74.623 60.504 74.707 ;
    END
  END Min_Wdata_ram[96]
  PIN Min_Wdata_ram[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.456 0 39.48 0.084 ;
    END
  END Min_Wdata_ram[97]
  PIN Min_Wdata_ram[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.968 0 55.992 0.084 ;
    END
  END Min_Wdata_ram[98]
  PIN Min_Wdata_ram[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.624 0 6.648 0.084 ;
    END
  END Min_Wdata_ram[99]
  PIN Min_Wdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.768 74.707 36.792 ;
    END
  END Min_Wdata_ram[9]
  PIN Min_addr_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.384 74.707 48.408 ;
    END
  END Min_addr_ram[0]
  PIN Min_addr_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.024 74.707 57.048 ;
    END
  END Min_addr_ram[10]
  PIN Min_addr_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.104 74.707 55.128 ;
    END
  END Min_addr_ram[11]
  PIN Min_addr_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.28 74.707 53.304 ;
    END
  END Min_addr_ram[12]
  PIN Min_addr_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.048 74.707 54.072 ;
    END
  END Min_addr_ram[13]
  PIN Min_addr_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.352 74.707 56.376 ;
    END
  END Min_addr_ram[14]
  PIN Min_addr_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.856 74.707 53.88 ;
    END
  END Min_addr_ram[15]
  PIN Min_addr_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.68 74.707 55.704 ;
    END
  END Min_addr_ram[16]
  PIN Min_addr_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.216 74.707 57.24 ;
    END
  END Min_addr_ram[17]
  PIN Min_addr_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.608 74.707 52.632 ;
    END
  END Min_addr_ram[18]
  PIN Min_addr_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.488 74.707 55.512 ;
    END
  END Min_addr_ram[19]
  PIN Min_addr_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.576 74.707 48.6 ;
    END
  END Min_addr_ram[1]
  PIN Min_addr_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.032 74.707 52.056 ;
    END
  END Min_addr_ram[20]
  PIN Min_addr_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.512 74.707 52.536 ;
    END
  END Min_addr_ram[21]
  PIN Min_addr_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.16 74.707 56.184 ;
    END
  END Min_addr_ram[22]
  PIN Min_addr_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.824 74.707 49.848 ;
    END
  END Min_addr_ram[23]
  PIN Min_addr_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.144 74.707 54.168 ;
    END
  END Min_addr_ram[24]
  PIN Min_addr_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.36 74.707 51.384 ;
    END
  END Min_addr_ram[25]
  PIN Min_addr_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.592 74.707 50.616 ;
    END
  END Min_addr_ram[26]
  PIN Min_addr_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.472 74.707 53.496 ;
    END
  END Min_addr_ram[27]
  PIN Min_addr_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.976 74.707 51 ;
    END
  END Min_addr_ram[28]
  PIN Min_addr_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.008 74.707 55.032 ;
    END
  END Min_addr_ram[29]
  PIN Min_addr_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.152 74.707 49.176 ;
    END
  END Min_addr_ram[2]
  PIN Min_addr_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.32 74.707 52.344 ;
    END
  END Min_addr_ram[30]
  PIN Min_addr_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.184 74.707 53.208 ;
    END
  END Min_addr_ram[31]
  PIN Min_addr_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.832 74.707 56.856 ;
    END
  END Min_addr_ram[32]
  PIN Min_addr_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.704 74.707 52.728 ;
    END
  END Min_addr_ram[33]
  PIN Min_addr_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.736 74.707 56.76 ;
    END
  END Min_addr_ram[34]
  PIN Min_addr_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.968 74.707 55.992 ;
    END
  END Min_addr_ram[35]
  PIN Min_addr_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.896 74.707 52.92 ;
    END
  END Min_addr_ram[36]
  PIN Min_addr_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.776 74.707 55.8 ;
    END
  END Min_addr_ram[37]
  PIN Min_addr_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.544 74.707 56.568 ;
    END
  END Min_addr_ram[38]
  PIN Min_addr_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.664 74.707 53.688 ;
    END
  END Min_addr_ram[39]
  PIN Min_addr_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.056 74.707 49.08 ;
    END
  END Min_addr_ram[3]
  PIN Min_addr_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.72 74.707 54.744 ;
    END
  END Min_addr_ram[40]
  PIN Min_addr_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.8 74.707 52.824 ;
    END
  END Min_addr_ram[41]
  PIN Min_addr_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.76 74.707 53.784 ;
    END
  END Min_addr_ram[42]
  PIN Min_addr_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.2 74.707 55.224 ;
    END
  END Min_addr_ram[43]
  PIN Min_addr_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.048 74.623 54.072 74.707 ;
    END
  END Min_addr_ram[44]
  PIN Min_addr_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.952 74.623 53.976 74.707 ;
    END
  END Min_addr_ram[45]
  PIN Min_addr_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.416 74.707 52.44 ;
    END
  END Min_addr_ram[4]
  PIN Min_addr_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.168 74.707 51.192 ;
    END
  END Min_addr_ram[5]
  PIN Min_addr_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.648 74.707 51.672 ;
    END
  END Min_addr_ram[6]
  PIN Min_addr_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.84 74.707 51.864 ;
    END
  END Min_addr_ram[7]
  PIN Min_addr_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.064 74.707 56.088 ;
    END
  END Min_addr_ram[8]
  PIN Min_addr_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.792 74.707 57.816 ;
    END
  END Min_addr_ram[9]
  PIN Min_data_ram_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.096 74.707 48.12 ;
    END
  END Min_data_ram_size[0]
  PIN Min_data_ram_size[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.96 74.707 48.984 ;
    END
  END Min_data_ram_size[10]
  PIN Min_data_ram_size[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.888 74.707 57.912 ;
    END
  END Min_data_ram_size[11]
  PIN Min_data_ram_size[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.504 74.707 57.528 ;
    END
  END Min_data_ram_size[12]
  PIN Min_data_ram_size[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.768 74.707 48.792 ;
    END
  END Min_data_ram_size[13]
  PIN Min_data_ram_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48 74.707 48.024 ;
    END
  END Min_data_ram_size[1]
  PIN Min_data_ram_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.904 74.707 47.928 ;
    END
  END Min_data_ram_size[2]
  PIN Min_data_ram_size[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.808 74.707 47.832 ;
    END
  END Min_data_ram_size[3]
  PIN Min_data_ram_size[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.632 74.707 49.656 ;
    END
  END Min_data_ram_size[4]
  PIN Min_data_ram_size[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.344 74.707 49.368 ;
    END
  END Min_data_ram_size[5]
  PIN Min_data_ram_size[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.728 74.707 49.752 ;
    END
  END Min_data_ram_size[6]
  PIN Min_data_ram_size[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.64 74.707 56.664 ;
    END
  END Min_data_ram_size[7]
  PIN Min_data_ram_size[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.392 74.707 55.416 ;
    END
  END Min_data_ram_size[8]
  PIN Min_data_ram_size[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.952 74.707 53.976 ;
    END
  END Min_data_ram_size[9]
  PIN Min_oe_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.712 74.707 47.736 ;
    END
  END Min_oe_ram[0]
  PIN Min_oe_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.192 74.707 48.216 ;
    END
  END Min_oe_ram[1]
  PIN Min_we_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.744 74.707 51.768 ;
    END
  END Min_we_ram[0]
  PIN Min_we_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  43.296 74.623 43.32 74.707 ;
    END
  END Min_we_ram[1]
  PIN Mout_Wdata_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.016 74.707 38.04 ;
    END
  END Mout_Wdata_ram[0]
  PIN Mout_Wdata_ram[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.664 74.623 53.688 74.707 ;
    END
  END Mout_Wdata_ram[100]
  PIN Mout_Wdata_ram[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.056 74.623 61.08 74.707 ;
    END
  END Mout_Wdata_ram[101]
  PIN Mout_Wdata_ram[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.744 0.084 3.768 ;
    END
  END Mout_Wdata_ram[102]
  PIN Mout_Wdata_ram[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.808 74.623 59.832 74.707 ;
    END
  END Mout_Wdata_ram[103]
  PIN Mout_Wdata_ram[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.728 74.623 13.752 74.707 ;
    END
  END Mout_Wdata_ram[104]
  PIN Mout_Wdata_ram[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.216 74.623 33.24 74.707 ;
    END
  END Mout_Wdata_ram[105]
  PIN Mout_Wdata_ram[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.272 0 58.296 0.084 ;
    END
  END Mout_Wdata_ram[106]
  PIN Mout_Wdata_ram[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.232 0 59.256 0.084 ;
    END
  END Mout_Wdata_ram[107]
  PIN Mout_Wdata_ram[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.816 74.623 6.84 74.707 ;
    END
  END Mout_Wdata_ram[108]
  PIN Mout_Wdata_ram[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.16 0 32.184 0.084 ;
    END
  END Mout_Wdata_ram[109]
  PIN Mout_Wdata_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.536 74.707 37.56 ;
    END
  END Mout_Wdata_ram[10]
  PIN Mout_Wdata_ram[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.048 0 54.072 0.084 ;
    END
  END Mout_Wdata_ram[110]
  PIN Mout_Wdata_ram[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.536 0 61.56 0.084 ;
    END
  END Mout_Wdata_ram[111]
  PIN Mout_Wdata_ram[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.592 0 62.616 0.084 ;
    END
  END Mout_Wdata_ram[112]
  PIN Mout_Wdata_ram[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 70.56 74.707 70.584 ;
    END
  END Mout_Wdata_ram[113]
  PIN Mout_Wdata_ram[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.368 74.623 34.392 74.707 ;
    END
  END Mout_Wdata_ram[114]
  PIN Mout_Wdata_ram[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.36 0 63.384 0.084 ;
    END
  END Mout_Wdata_ram[115]
  PIN Mout_Wdata_ram[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.52 74.623 59.544 74.707 ;
    END
  END Mout_Wdata_ram[116]
  PIN Mout_Wdata_ram[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.08 74.623 58.104 74.707 ;
    END
  END Mout_Wdata_ram[117]
  PIN Mout_Wdata_ram[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.112 74.623 38.136 74.707 ;
    END
  END Mout_Wdata_ram[118]
  PIN Mout_Wdata_ram[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.792 74.623 57.816 74.707 ;
    END
  END Mout_Wdata_ram[119]
  PIN Mout_Wdata_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.88 74.707 38.904 ;
    END
  END Mout_Wdata_ram[11]
  PIN Mout_Wdata_ram[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.88 0 62.904 0.084 ;
    END
  END Mout_Wdata_ram[120]
  PIN Mout_Wdata_ram[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.664 74.623 41.688 74.707 ;
    END
  END Mout_Wdata_ram[121]
  PIN Mout_Wdata_ram[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.36 0 39.384 0.084 ;
    END
  END Mout_Wdata_ram[122]
  PIN Mout_Wdata_ram[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.088 74.623 53.112 74.707 ;
    END
  END Mout_Wdata_ram[123]
  PIN Mout_Wdata_ram[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.632 0 61.656 0.084 ;
    END
  END Mout_Wdata_ram[124]
  PIN Mout_Wdata_ram[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.912 0 6.936 0.084 ;
    END
  END Mout_Wdata_ram[125]
  PIN Mout_Wdata_ram[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.768 0 36.792 0.084 ;
    END
  END Mout_Wdata_ram[126]
  PIN Mout_Wdata_ram[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.248 0 61.272 0.084 ;
    END
  END Mout_Wdata_ram[127]
  PIN Mout_Wdata_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 35.328 74.707 35.352 ;
    END
  END Mout_Wdata_ram[12]
  PIN Mout_Wdata_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.944 74.707 34.968 ;
    END
  END Mout_Wdata_ram[13]
  PIN Mout_Wdata_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.272 74.707 34.296 ;
    END
  END Mout_Wdata_ram[14]
  PIN Mout_Wdata_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.16 74.707 32.184 ;
    END
  END Mout_Wdata_ram[15]
  PIN Mout_Wdata_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.256 74.707 32.28 ;
    END
  END Mout_Wdata_ram[16]
  PIN Mout_Wdata_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.68 74.707 31.704 ;
    END
  END Mout_Wdata_ram[17]
  PIN Mout_Wdata_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.064 74.707 32.088 ;
    END
  END Mout_Wdata_ram[18]
  PIN Mout_Wdata_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.968 74.707 31.992 ;
    END
  END Mout_Wdata_ram[19]
  PIN Mout_Wdata_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.96 74.707 36.984 ;
    END
  END Mout_Wdata_ram[1]
  PIN Mout_Wdata_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.776 74.707 31.8 ;
    END
  END Mout_Wdata_ram[20]
  PIN Mout_Wdata_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.64 74.707 32.664 ;
    END
  END Mout_Wdata_ram[21]
  PIN Mout_Wdata_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 31.008 74.707 31.032 ;
    END
  END Mout_Wdata_ram[22]
  PIN Mout_Wdata_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.024 74.707 33.048 ;
    END
  END Mout_Wdata_ram[23]
  PIN Mout_Wdata_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 33.696 74.707 33.72 ;
    END
  END Mout_Wdata_ram[24]
  PIN Mout_Wdata_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 32.832 74.707 32.856 ;
    END
  END Mout_Wdata_ram[25]
  PIN Mout_Wdata_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.368 74.707 34.392 ;
    END
  END Mout_Wdata_ram[26]
  PIN Mout_Wdata_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 34.656 74.707 34.68 ;
    END
  END Mout_Wdata_ram[27]
  PIN Mout_Wdata_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.192 74.707 36.216 ;
    END
  END Mout_Wdata_ram[28]
  PIN Mout_Wdata_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.672 74.707 36.696 ;
    END
  END Mout_Wdata_ram[29]
  PIN Mout_Wdata_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.056 74.707 37.08 ;
    END
  END Mout_Wdata_ram[2]
  PIN Mout_Wdata_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.112 74.707 38.136 ;
    END
  END Mout_Wdata_ram[30]
  PIN Mout_Wdata_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.032 74.707 40.056 ;
    END
  END Mout_Wdata_ram[31]
  PIN Mout_Wdata_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.568 74.707 53.592 ;
    END
  END Mout_Wdata_ram[32]
  PIN Mout_Wdata_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  46.752 74.623 46.776 74.707 ;
    END
  END Mout_Wdata_ram[33]
  PIN Mout_Wdata_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.416 74.707 40.44 ;
    END
  END Mout_Wdata_ram[34]
  PIN Mout_Wdata_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.144 74.707 42.168 ;
    END
  END Mout_Wdata_ram[35]
  PIN Mout_Wdata_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.8 74.707 40.824 ;
    END
  END Mout_Wdata_ram[36]
  PIN Mout_Wdata_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 42.72 74.707 42.744 ;
    END
  END Mout_Wdata_ram[37]
  PIN Mout_Wdata_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.24 74.707 54.264 ;
    END
  END Mout_Wdata_ram[38]
  PIN Mout_Wdata_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.392 74.707 43.416 ;
    END
  END Mout_Wdata_ram[39]
  PIN Mout_Wdata_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.208 74.707 38.232 ;
    END
  END Mout_Wdata_ram[3]
  PIN Mout_Wdata_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.104 74.707 43.128 ;
    END
  END Mout_Wdata_ram[40]
  PIN Mout_Wdata_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.856 74.707 41.88 ;
    END
  END Mout_Wdata_ram[41]
  PIN Mout_Wdata_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.32 74.707 40.344 ;
    END
  END Mout_Wdata_ram[42]
  PIN Mout_Wdata_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.568 74.707 41.592 ;
    END
  END Mout_Wdata_ram[43]
  PIN Mout_Wdata_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.256 74.707 44.28 ;
    END
  END Mout_Wdata_ram[44]
  PIN Mout_Wdata_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.224 74.707 40.248 ;
    END
  END Mout_Wdata_ram[45]
  PIN Mout_Wdata_ram[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 47.616 74.707 47.64 ;
    END
  END Mout_Wdata_ram[46]
  PIN Mout_Wdata_ram[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.664 74.707 41.688 ;
    END
  END Mout_Wdata_ram[47]
  PIN Mout_Wdata_ram[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.872 74.707 43.896 ;
    END
  END Mout_Wdata_ram[48]
  PIN Mout_Wdata_ram[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.16 74.707 44.184 ;
    END
  END Mout_Wdata_ram[49]
  PIN Mout_Wdata_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 39.648 74.707 39.672 ;
    END
  END Mout_Wdata_ram[4]
  PIN Mout_Wdata_ram[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.608 74.707 40.632 ;
    END
  END Mout_Wdata_ram[50]
  PIN Mout_Wdata_ram[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.12 74.707 45.144 ;
    END
  END Mout_Wdata_ram[51]
  PIN Mout_Wdata_ram[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 41.952 74.707 41.976 ;
    END
  END Mout_Wdata_ram[52]
  PIN Mout_Wdata_ram[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.352 74.707 44.376 ;
    END
  END Mout_Wdata_ram[53]
  PIN Mout_Wdata_ram[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.296 74.707 43.32 ;
    END
  END Mout_Wdata_ram[54]
  PIN Mout_Wdata_ram[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.552 74.707 51.576 ;
    END
  END Mout_Wdata_ram[55]
  PIN Mout_Wdata_ram[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 46.944 74.707 46.968 ;
    END
  END Mout_Wdata_ram[56]
  PIN Mout_Wdata_ram[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.888 74.707 45.912 ;
    END
  END Mout_Wdata_ram[57]
  PIN Mout_Wdata_ram[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.696 74.707 45.72 ;
    END
  END Mout_Wdata_ram[58]
  PIN Mout_Wdata_ram[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.408 74.707 57.432 ;
    END
  END Mout_Wdata_ram[59]
  PIN Mout_Wdata_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.304 74.707 38.328 ;
    END
  END Mout_Wdata_ram[5]
  PIN Mout_Wdata_ram[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.408 74.707 45.432 ;
    END
  END Mout_Wdata_ram[60]
  PIN Mout_Wdata_ram[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 43.776 74.707 43.8 ;
    END
  END Mout_Wdata_ram[61]
  PIN Mout_Wdata_ram[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 44.832 74.707 44.856 ;
    END
  END Mout_Wdata_ram[62]
  PIN Mout_Wdata_ram[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 45.024 74.707 45.048 ;
    END
  END Mout_Wdata_ram[63]
  PIN Mout_Wdata_ram[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.136 74.623 23.16 74.707 ;
    END
  END Mout_Wdata_ram[64]
  PIN Mout_Wdata_ram[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.944 74.623 58.968 74.707 ;
    END
  END Mout_Wdata_ram[65]
  PIN Mout_Wdata_ram[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.848 74.623 58.872 74.707 ;
    END
  END Mout_Wdata_ram[66]
  PIN Mout_Wdata_ram[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  44.16 74.623 44.184 74.707 ;
    END
  END Mout_Wdata_ram[67]
  PIN Mout_Wdata_ram[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.752 0 34.776 0.084 ;
    END
  END Mout_Wdata_ram[68]
  PIN Mout_Wdata_ram[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.712 74.623 59.736 74.707 ;
    END
  END Mout_Wdata_ram[69]
  PIN Mout_Wdata_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 40.128 74.707 40.152 ;
    END
  END Mout_Wdata_ram[6]
  PIN Mout_Wdata_ram[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  66.72 74.623 66.744 74.707 ;
    END
  END Mout_Wdata_ram[70]
  PIN Mout_Wdata_ram[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  45.216 0 45.24 0.084 ;
    END
  END Mout_Wdata_ram[71]
  PIN Mout_Wdata_ram[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.576 74.623 60.6 74.707 ;
    END
  END Mout_Wdata_ram[72]
  PIN Mout_Wdata_ram[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.688 74.623 2.712 74.707 ;
    END
  END Mout_Wdata_ram[73]
  PIN Mout_Wdata_ram[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.472 74.623 53.496 74.707 ;
    END
  END Mout_Wdata_ram[74]
  PIN Mout_Wdata_ram[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.424 74.623 59.448 74.707 ;
    END
  END Mout_Wdata_ram[75]
  PIN Mout_Wdata_ram[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.28 0 17.304 0.084 ;
    END
  END Mout_Wdata_ram[76]
  PIN Mout_Wdata_ram[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.704 0 52.728 0.084 ;
    END
  END Mout_Wdata_ram[77]
  PIN Mout_Wdata_ram[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.896 74.623 52.92 74.707 ;
    END
  END Mout_Wdata_ram[78]
  PIN Mout_Wdata_ram[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.904 74.623 59.928 74.707 ;
    END
  END Mout_Wdata_ram[79]
  PIN Mout_Wdata_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.496 74.707 38.52 ;
    END
  END Mout_Wdata_ram[7]
  PIN Mout_Wdata_ram[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.72 74.623 54.744 74.707 ;
    END
  END Mout_Wdata_ram[80]
  PIN Mout_Wdata_ram[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.968 74.623 55.992 74.707 ;
    END
  END Mout_Wdata_ram[81]
  PIN Mout_Wdata_ram[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.656 0 34.68 0.084 ;
    END
  END Mout_Wdata_ram[82]
  PIN Mout_Wdata_ram[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.856 74.623 53.88 74.707 ;
    END
  END Mout_Wdata_ram[83]
  PIN Mout_Wdata_ram[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.576 0 60.6 0.084 ;
    END
  END Mout_Wdata_ram[84]
  PIN Mout_Wdata_ram[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.288 0 60.312 0.084 ;
    END
  END Mout_Wdata_ram[85]
  PIN Mout_Wdata_ram[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.408 74.623 21.432 74.707 ;
    END
  END Mout_Wdata_ram[86]
  PIN Mout_Wdata_ram[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  43.104 0 43.128 0.084 ;
    END
  END Mout_Wdata_ram[87]
  PIN Mout_Wdata_ram[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60 74.623 60.024 74.707 ;
    END
  END Mout_Wdata_ram[88]
  PIN Mout_Wdata_ram[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 62.784 74.707 62.808 ;
    END
  END Mout_Wdata_ram[89]
  PIN Mout_Wdata_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 37.824 74.707 37.848 ;
    END
  END Mout_Wdata_ram[8]
  PIN Mout_Wdata_ram[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  45.696 74.623 45.72 74.707 ;
    END
  END Mout_Wdata_ram[90]
  PIN Mout_Wdata_ram[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.376 74.623 41.4 74.707 ;
    END
  END Mout_Wdata_ram[91]
  PIN Mout_Wdata_ram[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.264 0 39.288 0.084 ;
    END
  END Mout_Wdata_ram[92]
  PIN Mout_Wdata_ram[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.552 0 63.576 0.084 ;
    END
  END Mout_Wdata_ram[93]
  PIN Mout_Wdata_ram[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.512 74.623 52.536 74.707 ;
    END
  END Mout_Wdata_ram[94]
  PIN Mout_Wdata_ram[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.272 74.623 58.296 74.707 ;
    END
  END Mout_Wdata_ram[95]
  PIN Mout_Wdata_ram[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.672 74.623 60.696 74.707 ;
    END
  END Mout_Wdata_ram[96]
  PIN Mout_Wdata_ram[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.648 0 39.672 0.084 ;
    END
  END Mout_Wdata_ram[97]
  PIN Mout_Wdata_ram[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  56.16 0 56.184 0.084 ;
    END
  END Mout_Wdata_ram[98]
  PIN Mout_Wdata_ram[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.816 0 6.84 0.084 ;
    END
  END Mout_Wdata_ram[99]
  PIN Mout_Wdata_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 36.864 74.707 36.888 ;
    END
  END Mout_Wdata_ram[9]
  PIN Mout_addr_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.672 74.707 48.696 ;
    END
  END Mout_addr_ram[0]
  PIN Mout_addr_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.376 74.707 53.4 ;
    END
  END Mout_addr_ram[10]
  PIN Mout_addr_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.928 74.707 56.952 ;
    END
  END Mout_addr_ram[11]
  PIN Mout_addr_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.872 74.707 55.896 ;
    END
  END Mout_addr_ram[12]
  PIN Mout_addr_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.624 74.707 54.648 ;
    END
  END Mout_addr_ram[13]
  PIN Mout_addr_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.528 74.707 54.552 ;
    END
  END Mout_addr_ram[14]
  PIN Mout_addr_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.296 74.707 55.32 ;
    END
  END Mout_addr_ram[15]
  PIN Mout_addr_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.696 74.707 57.72 ;
    END
  END Mout_addr_ram[16]
  PIN Mout_addr_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.312 74.707 57.336 ;
    END
  END Mout_addr_ram[17]
  PIN Mout_addr_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 53.088 74.707 53.112 ;
    END
  END Mout_addr_ram[18]
  PIN Mout_addr_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.336 74.707 54.36 ;
    END
  END Mout_addr_ram[19]
  PIN Mout_addr_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.016 74.707 50.04 ;
    END
  END Mout_addr_ram[1]
  PIN Mout_addr_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.936 74.707 51.96 ;
    END
  END Mout_addr_ram[20]
  PIN Mout_addr_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.08 74.707 58.104 ;
    END
  END Mout_addr_ram[21]
  PIN Mout_addr_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.176 74.707 58.2 ;
    END
  END Mout_addr_ram[22]
  PIN Mout_addr_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 57.6 74.707 57.624 ;
    END
  END Mout_addr_ram[23]
  PIN Mout_addr_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.864 74.707 48.888 ;
    END
  END Mout_addr_ram[24]
  PIN Mout_addr_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 49.44 74.707 49.464 ;
    END
  END Mout_addr_ram[25]
  PIN Mout_addr_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 50.784 74.707 50.808 ;
    END
  END Mout_addr_ram[26]
  PIN Mout_addr_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 52.992 74.707 53.016 ;
    END
  END Mout_addr_ram[27]
  PIN Mout_addr_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 51.072 74.707 51.096 ;
    END
  END Mout_addr_ram[28]
  PIN Mout_addr_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.432 74.707 54.456 ;
    END
  END Mout_addr_ram[29]
  PIN Mout_addr_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 48.48 74.707 48.504 ;
    END
  END Mout_addr_ram[2]
  PIN Mout_addr_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 56.256 74.707 56.28 ;
    END
  END Mout_addr_ram[30]
  PIN Mout_addr_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.816 74.707 54.84 ;
    END
  END Mout_addr_ram[31]
  PIN Mout_addr_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 54.912 74.707 54.936 ;
    END
  END Mout_addr_ram[32]
  PIN Mout_addr_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 55.584 74.707 55.608 ;
    END
  END Mout_addr_ram[33]
  PIN Mout_addr_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60.48 74.707 60.504 ;
    END
  END Mout_addr_ram[34]
  PIN Mout_addr_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  64.608 74.623 64.632 74.707 ;
    END
  END Mout_addr_ram[35]
  PIN Mout_addr_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.744 74.623 63.768 74.707 ;
    END
  END Mout_addr_ram[36]
  PIN Mout_addr_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.496 74.623 62.52 74.707 ;
    END
  END Mout_addr_ram[37]
  PIN Mout_addr_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.768 74.623 60.792 74.707 ;
    END
  END Mout_addr_ram[38]
  PIN Mout_addr_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  59.616 74.623 59.64 74.707 ;
    END
  END Mout_addr_ram[39]
  PIN Mout_addr_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.368 74.707 58.392 ;
    END
  END Mout_addr_ram[3]
  PIN Mout_addr_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.984 74.623 58.008 74.707 ;
    END
  END Mout_addr_ram[40]
  PIN Mout_addr_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.392 74.623 55.416 74.707 ;
    END
  END Mout_addr_ram[41]
  PIN Mout_addr_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.144 74.623 54.168 74.707 ;
    END
  END Mout_addr_ram[42]
  PIN Mout_addr_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  53.568 74.623 53.592 74.707 ;
    END
  END Mout_addr_ram[43]
  PIN Mout_addr_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.336 74.623 54.36 74.707 ;
    END
  END Mout_addr_ram[44]
  PIN Mout_addr_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.24 74.623 54.264 74.707 ;
    END
  END Mout_addr_ram[45]
  PIN Mout_addr_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.656 74.707 58.68 ;
    END
  END Mout_addr_ram[4]
  PIN Mout_addr_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.616 74.707 59.64 ;
    END
  END Mout_addr_ram[5]
  PIN Mout_addr_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60.192 74.707 60.216 ;
    END
  END Mout_addr_ram[6]
  PIN Mout_addr_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60.384 74.707 60.408 ;
    END
  END Mout_addr_ram[7]
  PIN Mout_addr_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.712 74.707 59.736 ;
    END
  END Mout_addr_ram[8]
  PIN Mout_addr_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.56 74.707 58.584 ;
    END
  END Mout_addr_ram[9]
  PIN Mout_data_ram_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.848 74.707 58.872 ;
    END
  END Mout_data_ram_size[0]
  PIN Mout_data_ram_size[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.104 74.623 55.128 74.707 ;
    END
  END Mout_data_ram_size[10]
  PIN Mout_data_ram_size[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.912 74.623 54.936 74.707 ;
    END
  END Mout_data_ram_size[11]
  PIN Mout_data_ram_size[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.816 74.623 54.84 74.707 ;
    END
  END Mout_data_ram_size[12]
  PIN Mout_data_ram_size[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.136 74.707 59.16 ;
    END
  END Mout_data_ram_size[13]
  PIN Mout_data_ram_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.808 74.707 59.832 ;
    END
  END Mout_data_ram_size[1]
  PIN Mout_data_ram_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.328 74.707 59.352 ;
    END
  END Mout_data_ram_size[2]
  PIN Mout_data_ram_size[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.944 74.707 58.968 ;
    END
  END Mout_data_ram_size[3]
  PIN Mout_data_ram_size[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.464 74.707 58.488 ;
    END
  END Mout_data_ram_size[4]
  PIN Mout_data_ram_size[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.272 74.707 58.296 ;
    END
  END Mout_data_ram_size[5]
  PIN Mout_data_ram_size[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  64.896 74.623 64.92 74.707 ;
    END
  END Mout_data_ram_size[6]
  PIN Mout_data_ram_size[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.008 74.623 55.032 74.707 ;
    END
  END Mout_data_ram_size[7]
  PIN Mout_data_ram_size[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.704 74.623 52.728 74.707 ;
    END
  END Mout_data_ram_size[8]
  PIN Mout_data_ram_size[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  52.8 74.623 52.824 74.707 ;
    END
  END Mout_data_ram_size[9]
  PIN Mout_oe_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.696 74.623 57.72 74.707 ;
    END
  END Mout_oe_ram[0]
  PIN Mout_oe_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.904 74.707 59.928 ;
    END
  END Mout_oe_ram[1]
  PIN Mout_we_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.784 74.707 38.808 ;
    END
  END Mout_we_ram[0]
  PIN Mout_we_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  43.488 74.623 43.512 74.707 ;
    END
  END Mout_we_ram[1]
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 64.992 0.084 65.016 ;
    END
  END clock
  PIN done_port
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.84 74.623 63.864 74.707 ;
    END
  END done_port
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.88 74.623 62.904 74.707 ;
    END
  END reset
  PIN start_port
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.92 74.623 61.944 74.707 ;
    END
  END start_port
  PIN vargs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  55.296 74.623 55.32 74.707 ;
    END
  END vargs[0]
  PIN vargs[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 58.752 74.707 58.776 ;
    END
  END vargs[10]
  PIN vargs[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  65.28 74.623 65.304 74.707 ;
    END
  END vargs[11]
  PIN vargs[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  64.704 74.623 64.728 74.707 ;
    END
  END vargs[12]
  PIN vargs[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  63.072 74.623 63.096 74.707 ;
    END
  END vargs[13]
  PIN vargs[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.112 74.623 62.136 74.707 ;
    END
  END vargs[14]
  PIN vargs[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.632 74.623 61.656 74.707 ;
    END
  END vargs[15]
  PIN vargs[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.176 74.623 58.2 74.707 ;
    END
  END vargs[16]
  PIN vargs[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.216 74.623 57.24 74.707 ;
    END
  END vargs[17]
  PIN vargs[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.024 74.623 57.048 74.707 ;
    END
  END vargs[18]
  PIN vargs[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.12 74.623 57.144 74.707 ;
    END
  END vargs[19]
  PIN vargs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.232 74.707 59.256 ;
    END
  END vargs[1]
  PIN vargs[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  56.928 74.623 56.952 74.707 ;
    END
  END vargs[20]
  PIN vargs[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  56.64 74.623 56.664 74.707 ;
    END
  END vargs[21]
  PIN vargs[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  56.736 74.623 56.76 74.707 ;
    END
  END vargs[22]
  PIN vargs[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.312 74.623 57.336 74.707 ;
    END
  END vargs[23]
  PIN vargs[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  57.408 74.623 57.432 74.707 ;
    END
  END vargs[24]
  PIN vargs[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.368 74.623 58.392 74.707 ;
    END
  END vargs[25]
  PIN vargs[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  58.464 74.623 58.488 74.707 ;
    END
  END vargs[26]
  PIN vargs[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  61.728 74.623 61.752 74.707 ;
    END
  END vargs[27]
  PIN vargs[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.96 74.623 60.984 74.707 ;
    END
  END vargs[28]
  PIN vargs[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.192 74.623 60.216 74.707 ;
    END
  END vargs[29]
  PIN vargs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 38.976 74.707 39 ;
    END
  END vargs[2]
  PIN vargs[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  60.384 74.623 60.408 74.707 ;
    END
  END vargs[30]
  PIN vargs[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.592 74.623 62.616 74.707 ;
    END
  END vargs[31]
  PIN vargs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  62.016 74.623 62.04 74.707 ;
    END
  END vargs[3]
  PIN vargs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60.288 74.707 60.312 ;
    END
  END vargs[4]
  PIN vargs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60 74.707 60.024 ;
    END
  END vargs[5]
  PIN vargs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.04 74.707 59.064 ;
    END
  END vargs[6]
  PIN vargs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.52 74.707 59.544 ;
    END
  END vargs[7]
  PIN vargs[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 59.424 74.707 59.448 ;
    END
  END vargs[8]
  PIN vargs[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  74.623 60.096 74.707 60.12 ;
    END
  END vargs[9]
  OBS
    LAYER M1 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M2 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M3 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M4 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M5 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M6 ;
     RECT  0 0 74.707 74.707 ;
    LAYER M7 ;
     RECT  0 0 74.707 74.707 ;
  END
END run_benchmark
END LIBRARY
