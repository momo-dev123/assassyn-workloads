VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA CSRFile_via1_2_28944_18_1_804_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 804 ;
END CSRFile_via1_2_28944_18_1_804_36_36

VIA CSRFile_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END CSRFile_VIA23_1_3_36_36

VIA CSRFile_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END CSRFile_VIA34_1_2_58_52

VIA CSRFile_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END CSRFile_VIA45_1_2_58_58

VIA CSRFile_via5_6_120_288_1_2_58_322
  VIARULE M6_M5widePWR1p152 ;
  CUTSIZE 0.024 0.288 ;
  LAYERS M5 V5 M6 ;
  CUTSPACING 0.034 0.034 ;
  ENCLOSURE 0.019 0 0 0 ;
  ROWCOL 1 2 ;
END CSRFile_via5_6_120_288_1_2_58_322

MACRO CSRFile
  FOREIGN CSRFile 0 0 ;
  CLASS BLOCK ;
  SIZE 31.005 BY 31.005 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.458 25.833 25.194 26.121 ;
        RECT  1.458 19.833 25.194 20.121 ;
        RECT  1.458 13.833 25.194 14.121 ;
        RECT  1.458 7.833 25.194 8.121 ;
        RECT  1.458 1.833 25.194 2.121 ;
      LAYER M5 ;
        RECT  25.074 1.327 25.194 29.993 ;
        RECT  19.17 1.327 19.29 29.993 ;
        RECT  13.266 1.327 13.386 29.993 ;
        RECT  7.362 1.327 7.482 29.993 ;
        RECT  1.458 1.327 1.578 29.993 ;
      LAYER M2 ;
        RECT  1.026 29.961 29.97 29.979 ;
        RECT  1.026 29.421 29.97 29.439 ;
        RECT  1.026 28.881 29.97 28.899 ;
        RECT  1.026 28.341 29.97 28.359 ;
        RECT  1.026 27.801 29.97 27.819 ;
        RECT  1.026 27.261 29.97 27.279 ;
        RECT  1.026 26.721 29.97 26.739 ;
        RECT  1.026 26.181 29.97 26.199 ;
        RECT  1.026 25.641 29.97 25.659 ;
        RECT  1.026 25.101 29.97 25.119 ;
        RECT  1.026 24.561 29.97 24.579 ;
        RECT  1.026 24.021 29.97 24.039 ;
        RECT  1.026 23.481 29.97 23.499 ;
        RECT  1.026 22.941 29.97 22.959 ;
        RECT  1.026 22.401 29.97 22.419 ;
        RECT  1.026 21.861 29.97 21.879 ;
        RECT  1.026 21.321 29.97 21.339 ;
        RECT  1.026 20.781 29.97 20.799 ;
        RECT  1.026 20.241 29.97 20.259 ;
        RECT  1.026 19.701 29.97 19.719 ;
        RECT  1.026 19.161 29.97 19.179 ;
        RECT  1.026 18.621 29.97 18.639 ;
        RECT  1.026 18.081 29.97 18.099 ;
        RECT  1.026 17.541 29.97 17.559 ;
        RECT  1.026 17.001 29.97 17.019 ;
        RECT  1.026 16.461 29.97 16.479 ;
        RECT  1.026 15.921 29.97 15.939 ;
        RECT  1.026 15.381 29.97 15.399 ;
        RECT  1.026 14.841 29.97 14.859 ;
        RECT  1.026 14.301 29.97 14.319 ;
        RECT  1.026 13.761 29.97 13.779 ;
        RECT  1.026 13.221 29.97 13.239 ;
        RECT  1.026 12.681 29.97 12.699 ;
        RECT  1.026 12.141 29.97 12.159 ;
        RECT  1.026 11.601 29.97 11.619 ;
        RECT  1.026 11.061 29.97 11.079 ;
        RECT  1.026 10.521 29.97 10.539 ;
        RECT  1.026 9.981 29.97 9.999 ;
        RECT  1.026 9.441 29.97 9.459 ;
        RECT  1.026 8.901 29.97 8.919 ;
        RECT  1.026 8.361 29.97 8.379 ;
        RECT  1.026 7.821 29.97 7.839 ;
        RECT  1.026 7.281 29.97 7.299 ;
        RECT  1.026 6.741 29.97 6.759 ;
        RECT  1.026 6.201 29.97 6.219 ;
        RECT  1.026 5.661 29.97 5.679 ;
        RECT  1.026 5.121 29.97 5.139 ;
        RECT  1.026 4.581 29.97 4.599 ;
        RECT  1.026 4.041 29.97 4.059 ;
        RECT  1.026 3.501 29.97 3.519 ;
        RECT  1.026 2.961 29.97 2.979 ;
        RECT  1.026 2.421 29.97 2.439 ;
        RECT  1.026 1.881 29.97 1.899 ;
        RECT  1.026 1.341 29.97 1.359 ;
      LAYER M1 ;
        RECT  1.026 29.961 29.97 29.979 ;
        RECT  1.026 29.421 29.97 29.439 ;
        RECT  1.026 28.881 29.97 28.899 ;
        RECT  1.026 28.341 29.97 28.359 ;
        RECT  1.026 27.801 29.97 27.819 ;
        RECT  1.026 27.261 29.97 27.279 ;
        RECT  1.026 26.721 29.97 26.739 ;
        RECT  1.026 26.181 29.97 26.199 ;
        RECT  1.026 25.641 29.97 25.659 ;
        RECT  1.026 25.101 29.97 25.119 ;
        RECT  1.026 24.561 29.97 24.579 ;
        RECT  1.026 24.021 29.97 24.039 ;
        RECT  1.026 23.481 29.97 23.499 ;
        RECT  1.026 22.941 29.97 22.959 ;
        RECT  1.026 22.401 29.97 22.419 ;
        RECT  1.026 21.861 29.97 21.879 ;
        RECT  1.026 21.321 29.97 21.339 ;
        RECT  1.026 20.781 29.97 20.799 ;
        RECT  1.026 20.241 29.97 20.259 ;
        RECT  1.026 19.701 29.97 19.719 ;
        RECT  1.026 19.161 29.97 19.179 ;
        RECT  1.026 18.621 29.97 18.639 ;
        RECT  1.026 18.081 29.97 18.099 ;
        RECT  1.026 17.541 29.97 17.559 ;
        RECT  1.026 17.001 29.97 17.019 ;
        RECT  1.026 16.461 29.97 16.479 ;
        RECT  1.026 15.921 29.97 15.939 ;
        RECT  1.026 15.381 29.97 15.399 ;
        RECT  1.026 14.841 29.97 14.859 ;
        RECT  1.026 14.301 29.97 14.319 ;
        RECT  1.026 13.761 29.97 13.779 ;
        RECT  1.026 13.221 29.97 13.239 ;
        RECT  1.026 12.681 29.97 12.699 ;
        RECT  1.026 12.141 29.97 12.159 ;
        RECT  1.026 11.601 29.97 11.619 ;
        RECT  1.026 11.061 29.97 11.079 ;
        RECT  1.026 10.521 29.97 10.539 ;
        RECT  1.026 9.981 29.97 9.999 ;
        RECT  1.026 9.441 29.97 9.459 ;
        RECT  1.026 8.901 29.97 8.919 ;
        RECT  1.026 8.361 29.97 8.379 ;
        RECT  1.026 7.821 29.97 7.839 ;
        RECT  1.026 7.281 29.97 7.299 ;
        RECT  1.026 6.741 29.97 6.759 ;
        RECT  1.026 6.201 29.97 6.219 ;
        RECT  1.026 5.661 29.97 5.679 ;
        RECT  1.026 5.121 29.97 5.139 ;
        RECT  1.026 4.581 29.97 4.599 ;
        RECT  1.026 4.041 29.97 4.059 ;
        RECT  1.026 3.501 29.97 3.519 ;
        RECT  1.026 2.961 29.97 2.979 ;
        RECT  1.026 2.421 29.97 2.439 ;
        RECT  1.026 1.881 29.97 1.899 ;
        RECT  1.026 1.341 29.97 1.359 ;
      VIA 25.134 25.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 19.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 13.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 7.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 1.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 25.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 19.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 13.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 7.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 1.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 25.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 19.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 13.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 7.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 1.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 25.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 19.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 13.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 7.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 1.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 25.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 19.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 13.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 7.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 1.977 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 29.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.953 25.179 29.987 ;
      VIA 25.134 29.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 29.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 29.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.413 25.179 29.447 ;
      VIA 25.134 29.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 29.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 28.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.873 25.179 28.907 ;
      VIA 25.134 28.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 28.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 28.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.333 25.179 28.367 ;
      VIA 25.134 28.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 28.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 27.81 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.793 25.179 27.827 ;
      VIA 25.134 27.81 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 27.81 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 27.27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.253 25.179 27.287 ;
      VIA 25.134 27.27 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 27.27 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 26.73 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.713 25.179 26.747 ;
      VIA 25.134 26.73 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 26.73 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 26.19 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.173 25.179 26.207 ;
      VIA 25.134 26.19 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 26.19 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 25.65 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.633 25.179 25.667 ;
      VIA 25.134 25.65 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 25.65 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 25.11 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.093 25.179 25.127 ;
      VIA 25.134 25.11 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 25.11 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 24.57 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.553 25.179 24.587 ;
      VIA 25.134 24.57 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 24.57 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 24.03 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.013 25.179 24.047 ;
      VIA 25.134 24.03 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 24.03 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 23.49 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 23.473 25.179 23.507 ;
      VIA 25.134 23.49 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 23.49 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 22.95 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.933 25.179 22.967 ;
      VIA 25.134 22.95 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 22.95 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 22.41 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.393 25.179 22.427 ;
      VIA 25.134 22.41 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 22.41 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 21.87 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.853 25.179 21.887 ;
      VIA 25.134 21.87 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 21.87 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 21.33 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.313 25.179 21.347 ;
      VIA 25.134 21.33 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 21.33 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 20.79 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.773 25.179 20.807 ;
      VIA 25.134 20.79 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 20.79 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 20.25 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.233 25.179 20.267 ;
      VIA 25.134 20.25 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 20.25 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 19.71 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.693 25.179 19.727 ;
      VIA 25.134 19.71 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 19.71 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 19.17 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.153 25.179 19.187 ;
      VIA 25.134 19.17 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 19.17 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 18.63 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.613 25.179 18.647 ;
      VIA 25.134 18.63 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 18.63 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 18.09 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.073 25.179 18.107 ;
      VIA 25.134 18.09 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 18.09 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 17.55 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 17.533 25.179 17.567 ;
      VIA 25.134 17.55 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 17.55 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 17.01 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.993 25.179 17.027 ;
      VIA 25.134 17.01 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 17.01 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 16.47 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.453 25.179 16.487 ;
      VIA 25.134 16.47 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 16.47 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 15.93 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.913 25.179 15.947 ;
      VIA 25.134 15.93 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 15.93 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 15.39 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.373 25.179 15.407 ;
      VIA 25.134 15.39 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 15.39 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 14.85 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.833 25.179 14.867 ;
      VIA 25.134 14.85 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 14.85 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 14.31 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.293 25.179 14.327 ;
      VIA 25.134 14.31 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 14.31 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 13.77 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.753 25.179 13.787 ;
      VIA 25.134 13.77 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 13.77 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 13.23 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.213 25.179 13.247 ;
      VIA 25.134 13.23 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 13.23 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 12.69 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.673 25.179 12.707 ;
      VIA 25.134 12.69 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 12.69 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 12.15 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.133 25.179 12.167 ;
      VIA 25.134 12.15 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 12.15 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 11.61 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.593 25.179 11.627 ;
      VIA 25.134 11.61 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 11.61 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 11.07 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.053 25.179 11.087 ;
      VIA 25.134 11.07 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 11.07 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 10.53 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 10.513 25.179 10.547 ;
      VIA 25.134 10.53 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 10.53 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 9.99 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.973 25.179 10.007 ;
      VIA 25.134 9.99 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 9.99 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 9.45 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.433 25.179 9.467 ;
      VIA 25.134 9.45 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 9.45 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 8.91 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.893 25.179 8.927 ;
      VIA 25.134 8.91 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 8.91 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 8.37 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.353 25.179 8.387 ;
      VIA 25.134 8.37 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 8.37 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 7.83 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.813 25.179 7.847 ;
      VIA 25.134 7.83 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 7.83 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 7.29 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.273 25.179 7.307 ;
      VIA 25.134 7.29 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 7.29 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 6.75 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.733 25.179 6.767 ;
      VIA 25.134 6.75 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 6.75 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 6.21 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.193 25.179 6.227 ;
      VIA 25.134 6.21 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 6.21 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 5.67 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.653 25.179 5.687 ;
      VIA 25.134 5.67 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 5.67 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 5.13 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.113 25.179 5.147 ;
      VIA 25.134 5.13 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 5.13 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 4.59 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.573 25.179 4.607 ;
      VIA 25.134 4.59 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 4.59 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 4.05 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.033 25.179 4.067 ;
      VIA 25.134 4.05 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 4.05 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 3.51 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 3.493 25.179 3.527 ;
      VIA 25.134 3.51 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 3.51 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 2.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.953 25.179 2.987 ;
      VIA 25.134 2.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 2.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 2.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.413 25.179 2.447 ;
      VIA 25.134 2.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 2.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 1.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.873 25.179 1.907 ;
      VIA 25.134 1.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 1.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 25.134 1.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.333 25.179 1.367 ;
      VIA 25.134 1.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 25.134 1.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 29.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.953 19.275 29.987 ;
      VIA 19.23 29.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 29.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 29.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.413 19.275 29.447 ;
      VIA 19.23 29.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 29.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 28.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.873 19.275 28.907 ;
      VIA 19.23 28.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 28.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 28.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.333 19.275 28.367 ;
      VIA 19.23 28.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 28.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 27.81 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.793 19.275 27.827 ;
      VIA 19.23 27.81 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 27.81 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 27.27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.253 19.275 27.287 ;
      VIA 19.23 27.27 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 27.27 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 26.73 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.713 19.275 26.747 ;
      VIA 19.23 26.73 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 26.73 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 26.19 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.173 19.275 26.207 ;
      VIA 19.23 26.19 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 26.19 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 25.65 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.633 19.275 25.667 ;
      VIA 19.23 25.65 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 25.65 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 25.11 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.093 19.275 25.127 ;
      VIA 19.23 25.11 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 25.11 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 24.57 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.553 19.275 24.587 ;
      VIA 19.23 24.57 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 24.57 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 24.03 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.013 19.275 24.047 ;
      VIA 19.23 24.03 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 24.03 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 23.49 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 23.473 19.275 23.507 ;
      VIA 19.23 23.49 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 23.49 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 22.95 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.933 19.275 22.967 ;
      VIA 19.23 22.95 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 22.95 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 22.41 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.393 19.275 22.427 ;
      VIA 19.23 22.41 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 22.41 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 21.87 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.853 19.275 21.887 ;
      VIA 19.23 21.87 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 21.87 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 21.33 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.313 19.275 21.347 ;
      VIA 19.23 21.33 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 21.33 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 20.79 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.773 19.275 20.807 ;
      VIA 19.23 20.79 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 20.79 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 20.25 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.233 19.275 20.267 ;
      VIA 19.23 20.25 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 20.25 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 19.71 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.693 19.275 19.727 ;
      VIA 19.23 19.71 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 19.71 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 19.17 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.153 19.275 19.187 ;
      VIA 19.23 19.17 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 19.17 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 18.63 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.613 19.275 18.647 ;
      VIA 19.23 18.63 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 18.63 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 18.09 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.073 19.275 18.107 ;
      VIA 19.23 18.09 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 18.09 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 17.55 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 17.533 19.275 17.567 ;
      VIA 19.23 17.55 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 17.55 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 17.01 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.993 19.275 17.027 ;
      VIA 19.23 17.01 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 17.01 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 16.47 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.453 19.275 16.487 ;
      VIA 19.23 16.47 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 16.47 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 15.93 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.913 19.275 15.947 ;
      VIA 19.23 15.93 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 15.93 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 15.39 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.373 19.275 15.407 ;
      VIA 19.23 15.39 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 15.39 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 14.85 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.833 19.275 14.867 ;
      VIA 19.23 14.85 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 14.85 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 14.31 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.293 19.275 14.327 ;
      VIA 19.23 14.31 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 14.31 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 13.77 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.753 19.275 13.787 ;
      VIA 19.23 13.77 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 13.77 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 13.23 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.213 19.275 13.247 ;
      VIA 19.23 13.23 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 13.23 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 12.69 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.673 19.275 12.707 ;
      VIA 19.23 12.69 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 12.69 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 12.15 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.133 19.275 12.167 ;
      VIA 19.23 12.15 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 12.15 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 11.61 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.593 19.275 11.627 ;
      VIA 19.23 11.61 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 11.61 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 11.07 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.053 19.275 11.087 ;
      VIA 19.23 11.07 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 11.07 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 10.53 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 10.513 19.275 10.547 ;
      VIA 19.23 10.53 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 10.53 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 9.99 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.973 19.275 10.007 ;
      VIA 19.23 9.99 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 9.99 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 9.45 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.433 19.275 9.467 ;
      VIA 19.23 9.45 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 9.45 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 8.91 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.893 19.275 8.927 ;
      VIA 19.23 8.91 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 8.91 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 8.37 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.353 19.275 8.387 ;
      VIA 19.23 8.37 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 8.37 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 7.83 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.813 19.275 7.847 ;
      VIA 19.23 7.83 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 7.83 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 7.29 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.273 19.275 7.307 ;
      VIA 19.23 7.29 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 7.29 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 6.75 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.733 19.275 6.767 ;
      VIA 19.23 6.75 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 6.75 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 6.21 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.193 19.275 6.227 ;
      VIA 19.23 6.21 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 6.21 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 5.67 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.653 19.275 5.687 ;
      VIA 19.23 5.67 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 5.67 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 5.13 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.113 19.275 5.147 ;
      VIA 19.23 5.13 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 5.13 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 4.59 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.573 19.275 4.607 ;
      VIA 19.23 4.59 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 4.59 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 4.05 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.033 19.275 4.067 ;
      VIA 19.23 4.05 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 4.05 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 3.51 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 3.493 19.275 3.527 ;
      VIA 19.23 3.51 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 3.51 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 2.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.953 19.275 2.987 ;
      VIA 19.23 2.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 2.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 2.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.413 19.275 2.447 ;
      VIA 19.23 2.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 2.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 1.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.873 19.275 1.907 ;
      VIA 19.23 1.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 1.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.23 1.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.333 19.275 1.367 ;
      VIA 19.23 1.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.23 1.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 29.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.953 13.371 29.987 ;
      VIA 13.326 29.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 29.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 29.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.413 13.371 29.447 ;
      VIA 13.326 29.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 29.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 28.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.873 13.371 28.907 ;
      VIA 13.326 28.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 28.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 28.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.333 13.371 28.367 ;
      VIA 13.326 28.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 28.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 27.81 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.793 13.371 27.827 ;
      VIA 13.326 27.81 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 27.81 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 27.27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.253 13.371 27.287 ;
      VIA 13.326 27.27 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 27.27 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 26.73 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.713 13.371 26.747 ;
      VIA 13.326 26.73 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 26.73 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 26.19 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.173 13.371 26.207 ;
      VIA 13.326 26.19 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 26.19 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 25.65 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.633 13.371 25.667 ;
      VIA 13.326 25.65 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 25.65 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 25.11 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.093 13.371 25.127 ;
      VIA 13.326 25.11 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 25.11 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 24.57 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.553 13.371 24.587 ;
      VIA 13.326 24.57 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 24.57 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 24.03 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.013 13.371 24.047 ;
      VIA 13.326 24.03 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 24.03 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 23.49 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 23.473 13.371 23.507 ;
      VIA 13.326 23.49 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 23.49 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 22.95 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.933 13.371 22.967 ;
      VIA 13.326 22.95 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 22.95 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 22.41 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.393 13.371 22.427 ;
      VIA 13.326 22.41 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 22.41 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 21.87 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.853 13.371 21.887 ;
      VIA 13.326 21.87 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 21.87 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 21.33 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.313 13.371 21.347 ;
      VIA 13.326 21.33 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 21.33 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 20.79 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.773 13.371 20.807 ;
      VIA 13.326 20.79 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 20.79 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 20.25 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.233 13.371 20.267 ;
      VIA 13.326 20.25 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 20.25 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 19.71 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.693 13.371 19.727 ;
      VIA 13.326 19.71 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 19.71 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 19.17 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.153 13.371 19.187 ;
      VIA 13.326 19.17 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 19.17 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 18.63 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.613 13.371 18.647 ;
      VIA 13.326 18.63 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 18.63 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 18.09 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.073 13.371 18.107 ;
      VIA 13.326 18.09 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 18.09 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 17.55 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 17.533 13.371 17.567 ;
      VIA 13.326 17.55 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 17.55 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 17.01 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.993 13.371 17.027 ;
      VIA 13.326 17.01 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 17.01 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 16.47 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.453 13.371 16.487 ;
      VIA 13.326 16.47 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 16.47 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 15.93 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.913 13.371 15.947 ;
      VIA 13.326 15.93 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 15.93 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 15.39 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.373 13.371 15.407 ;
      VIA 13.326 15.39 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 15.39 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 14.85 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.833 13.371 14.867 ;
      VIA 13.326 14.85 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 14.85 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 14.31 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.293 13.371 14.327 ;
      VIA 13.326 14.31 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 14.31 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 13.77 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.753 13.371 13.787 ;
      VIA 13.326 13.77 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 13.77 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 13.23 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.213 13.371 13.247 ;
      VIA 13.326 13.23 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 13.23 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 12.69 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.673 13.371 12.707 ;
      VIA 13.326 12.69 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 12.69 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 12.15 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.133 13.371 12.167 ;
      VIA 13.326 12.15 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 12.15 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 11.61 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.593 13.371 11.627 ;
      VIA 13.326 11.61 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 11.61 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 11.07 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.053 13.371 11.087 ;
      VIA 13.326 11.07 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 11.07 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 10.53 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 10.513 13.371 10.547 ;
      VIA 13.326 10.53 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 10.53 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 9.99 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.973 13.371 10.007 ;
      VIA 13.326 9.99 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 9.99 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 9.45 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.433 13.371 9.467 ;
      VIA 13.326 9.45 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 9.45 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 8.91 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.893 13.371 8.927 ;
      VIA 13.326 8.91 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 8.91 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 8.37 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.353 13.371 8.387 ;
      VIA 13.326 8.37 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 8.37 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 7.83 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.813 13.371 7.847 ;
      VIA 13.326 7.83 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 7.83 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 7.29 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.273 13.371 7.307 ;
      VIA 13.326 7.29 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 7.29 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 6.75 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.733 13.371 6.767 ;
      VIA 13.326 6.75 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 6.75 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 6.21 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.193 13.371 6.227 ;
      VIA 13.326 6.21 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 6.21 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 5.67 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.653 13.371 5.687 ;
      VIA 13.326 5.67 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 5.67 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 5.13 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.113 13.371 5.147 ;
      VIA 13.326 5.13 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 5.13 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 4.59 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.573 13.371 4.607 ;
      VIA 13.326 4.59 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 4.59 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 4.05 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.033 13.371 4.067 ;
      VIA 13.326 4.05 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 4.05 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 3.51 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 3.493 13.371 3.527 ;
      VIA 13.326 3.51 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 3.51 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 2.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.953 13.371 2.987 ;
      VIA 13.326 2.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 2.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 2.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.413 13.371 2.447 ;
      VIA 13.326 2.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 2.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 1.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.873 13.371 1.907 ;
      VIA 13.326 1.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 1.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.326 1.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.333 13.371 1.367 ;
      VIA 13.326 1.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.326 1.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 29.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.953 7.467 29.987 ;
      VIA 7.422 29.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 29.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 29.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.413 7.467 29.447 ;
      VIA 7.422 29.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 29.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 28.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.873 7.467 28.907 ;
      VIA 7.422 28.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 28.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 28.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.333 7.467 28.367 ;
      VIA 7.422 28.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 28.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 27.81 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.793 7.467 27.827 ;
      VIA 7.422 27.81 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 27.81 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 27.27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.253 7.467 27.287 ;
      VIA 7.422 27.27 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 27.27 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 26.73 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.713 7.467 26.747 ;
      VIA 7.422 26.73 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 26.73 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 26.19 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.173 7.467 26.207 ;
      VIA 7.422 26.19 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 26.19 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 25.65 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.633 7.467 25.667 ;
      VIA 7.422 25.65 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 25.65 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 25.11 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.093 7.467 25.127 ;
      VIA 7.422 25.11 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 25.11 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 24.57 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.553 7.467 24.587 ;
      VIA 7.422 24.57 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 24.57 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 24.03 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.013 7.467 24.047 ;
      VIA 7.422 24.03 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 24.03 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 23.49 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 23.473 7.467 23.507 ;
      VIA 7.422 23.49 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 23.49 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 22.95 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.933 7.467 22.967 ;
      VIA 7.422 22.95 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 22.95 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 22.41 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.393 7.467 22.427 ;
      VIA 7.422 22.41 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 22.41 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 21.87 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.853 7.467 21.887 ;
      VIA 7.422 21.87 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 21.87 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 21.33 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.313 7.467 21.347 ;
      VIA 7.422 21.33 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 21.33 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 20.79 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.773 7.467 20.807 ;
      VIA 7.422 20.79 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 20.79 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 20.25 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.233 7.467 20.267 ;
      VIA 7.422 20.25 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 20.25 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 19.71 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.693 7.467 19.727 ;
      VIA 7.422 19.71 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 19.71 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 19.17 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.153 7.467 19.187 ;
      VIA 7.422 19.17 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 19.17 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 18.63 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.613 7.467 18.647 ;
      VIA 7.422 18.63 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 18.63 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 18.09 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.073 7.467 18.107 ;
      VIA 7.422 18.09 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 18.09 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 17.55 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 17.533 7.467 17.567 ;
      VIA 7.422 17.55 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 17.55 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 17.01 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.993 7.467 17.027 ;
      VIA 7.422 17.01 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 17.01 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 16.47 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.453 7.467 16.487 ;
      VIA 7.422 16.47 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 16.47 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 15.93 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.913 7.467 15.947 ;
      VIA 7.422 15.93 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 15.93 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 15.39 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.373 7.467 15.407 ;
      VIA 7.422 15.39 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 15.39 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 14.85 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.833 7.467 14.867 ;
      VIA 7.422 14.85 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 14.85 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 14.31 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.293 7.467 14.327 ;
      VIA 7.422 14.31 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 14.31 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 13.77 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.753 7.467 13.787 ;
      VIA 7.422 13.77 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 13.77 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 13.23 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.213 7.467 13.247 ;
      VIA 7.422 13.23 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 13.23 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 12.69 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.673 7.467 12.707 ;
      VIA 7.422 12.69 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 12.69 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 12.15 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.133 7.467 12.167 ;
      VIA 7.422 12.15 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 12.15 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 11.61 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.593 7.467 11.627 ;
      VIA 7.422 11.61 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 11.61 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 11.07 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.053 7.467 11.087 ;
      VIA 7.422 11.07 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 11.07 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 10.53 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 10.513 7.467 10.547 ;
      VIA 7.422 10.53 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 10.53 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 9.99 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.973 7.467 10.007 ;
      VIA 7.422 9.99 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 9.99 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 9.45 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.433 7.467 9.467 ;
      VIA 7.422 9.45 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 9.45 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 8.91 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.893 7.467 8.927 ;
      VIA 7.422 8.91 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 8.91 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 8.37 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.353 7.467 8.387 ;
      VIA 7.422 8.37 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 8.37 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 7.83 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.813 7.467 7.847 ;
      VIA 7.422 7.83 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 7.83 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 7.29 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.273 7.467 7.307 ;
      VIA 7.422 7.29 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 7.29 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 6.75 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.733 7.467 6.767 ;
      VIA 7.422 6.75 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 6.75 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 6.21 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.193 7.467 6.227 ;
      VIA 7.422 6.21 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 6.21 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 5.67 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.653 7.467 5.687 ;
      VIA 7.422 5.67 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 5.67 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 5.13 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.113 7.467 5.147 ;
      VIA 7.422 5.13 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 5.13 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 4.59 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.573 7.467 4.607 ;
      VIA 7.422 4.59 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 4.59 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 4.05 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.033 7.467 4.067 ;
      VIA 7.422 4.05 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 4.05 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 3.51 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 3.493 7.467 3.527 ;
      VIA 7.422 3.51 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 3.51 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 2.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.953 7.467 2.987 ;
      VIA 7.422 2.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 2.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 2.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.413 7.467 2.447 ;
      VIA 7.422 2.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 2.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 1.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.873 7.467 1.907 ;
      VIA 7.422 1.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 1.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.422 1.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.333 7.467 1.367 ;
      VIA 7.422 1.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.422 1.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 29.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.953 1.563 29.987 ;
      VIA 1.518 29.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 29.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 29.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.413 1.563 29.447 ;
      VIA 1.518 29.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 29.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 28.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.873 1.563 28.907 ;
      VIA 1.518 28.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 28.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 28.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.333 1.563 28.367 ;
      VIA 1.518 28.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 28.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 27.81 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.793 1.563 27.827 ;
      VIA 1.518 27.81 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 27.81 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 27.27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.253 1.563 27.287 ;
      VIA 1.518 27.27 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 27.27 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 26.73 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.713 1.563 26.747 ;
      VIA 1.518 26.73 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 26.73 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 26.19 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.173 1.563 26.207 ;
      VIA 1.518 26.19 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 26.19 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 25.65 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.633 1.563 25.667 ;
      VIA 1.518 25.65 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 25.65 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 25.11 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.093 1.563 25.127 ;
      VIA 1.518 25.11 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 25.11 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 24.57 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.553 1.563 24.587 ;
      VIA 1.518 24.57 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 24.57 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 24.03 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.013 1.563 24.047 ;
      VIA 1.518 24.03 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 24.03 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 23.49 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 23.473 1.563 23.507 ;
      VIA 1.518 23.49 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 23.49 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 22.95 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.933 1.563 22.967 ;
      VIA 1.518 22.95 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 22.95 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 22.41 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.393 1.563 22.427 ;
      VIA 1.518 22.41 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 22.41 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 21.87 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.853 1.563 21.887 ;
      VIA 1.518 21.87 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 21.87 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 21.33 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.313 1.563 21.347 ;
      VIA 1.518 21.33 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 21.33 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 20.79 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.773 1.563 20.807 ;
      VIA 1.518 20.79 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 20.79 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 20.25 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.233 1.563 20.267 ;
      VIA 1.518 20.25 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 20.25 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 19.71 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.693 1.563 19.727 ;
      VIA 1.518 19.71 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 19.71 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 19.17 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.153 1.563 19.187 ;
      VIA 1.518 19.17 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 19.17 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 18.63 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.613 1.563 18.647 ;
      VIA 1.518 18.63 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 18.63 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 18.09 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.073 1.563 18.107 ;
      VIA 1.518 18.09 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 18.09 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 17.55 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 17.533 1.563 17.567 ;
      VIA 1.518 17.55 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 17.55 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 17.01 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.993 1.563 17.027 ;
      VIA 1.518 17.01 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 17.01 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 16.47 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.453 1.563 16.487 ;
      VIA 1.518 16.47 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 16.47 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 15.93 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.913 1.563 15.947 ;
      VIA 1.518 15.93 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 15.93 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 15.39 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.373 1.563 15.407 ;
      VIA 1.518 15.39 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 15.39 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 14.85 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.833 1.563 14.867 ;
      VIA 1.518 14.85 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 14.85 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 14.31 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.293 1.563 14.327 ;
      VIA 1.518 14.31 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 14.31 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 13.77 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.753 1.563 13.787 ;
      VIA 1.518 13.77 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 13.77 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 13.23 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.213 1.563 13.247 ;
      VIA 1.518 13.23 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 13.23 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 12.69 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.673 1.563 12.707 ;
      VIA 1.518 12.69 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 12.69 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 12.15 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.133 1.563 12.167 ;
      VIA 1.518 12.15 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 12.15 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 11.61 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.593 1.563 11.627 ;
      VIA 1.518 11.61 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 11.61 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 11.07 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.053 1.563 11.087 ;
      VIA 1.518 11.07 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 11.07 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 10.53 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 10.513 1.563 10.547 ;
      VIA 1.518 10.53 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 10.53 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 9.99 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.973 1.563 10.007 ;
      VIA 1.518 9.99 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 9.99 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 9.45 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.433 1.563 9.467 ;
      VIA 1.518 9.45 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 9.45 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 8.91 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.893 1.563 8.927 ;
      VIA 1.518 8.91 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 8.91 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 8.37 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.353 1.563 8.387 ;
      VIA 1.518 8.37 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 8.37 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 7.83 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.813 1.563 7.847 ;
      VIA 1.518 7.83 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 7.83 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 7.29 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.273 1.563 7.307 ;
      VIA 1.518 7.29 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 7.29 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 6.75 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.733 1.563 6.767 ;
      VIA 1.518 6.75 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 6.75 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 6.21 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.193 1.563 6.227 ;
      VIA 1.518 6.21 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 6.21 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 5.67 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.653 1.563 5.687 ;
      VIA 1.518 5.67 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 5.67 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 5.13 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.113 1.563 5.147 ;
      VIA 1.518 5.13 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 5.13 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 4.59 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 CSRFile_VIA23_1_3_36_36 ;
      VIA 15.498 29.97 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 29.43 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 28.89 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 28.35 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 27.81 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 27.27 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 26.73 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 26.19 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 25.65 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 25.11 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 24.57 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 24.03 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 23.49 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 22.95 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 22.41 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 21.87 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 21.33 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 20.79 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 20.25 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 19.71 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 19.17 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 18.63 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 18.09 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 17.55 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 17.01 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 16.47 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 15.93 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 15.39 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 14.85 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 14.31 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 13.77 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 13.23 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 12.69 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 12.15 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 11.61 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 11.07 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 10.53 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 9.99 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 9.45 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 8.91 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 8.37 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 7.83 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 7.29 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 6.75 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 6.21 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 5.67 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 5.13 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 4.59 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 4.05 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 3.51 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 2.97 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 2.43 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 1.89 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 1.35 CSRFile_via1_2_28944_18_1_804_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.266 25.449 25.002 25.737 ;
        RECT  1.266 19.449 25.002 19.737 ;
        RECT  1.266 13.449 25.002 13.737 ;
        RECT  1.266 7.449 25.002 7.737 ;
        RECT  1.266 1.449 25.002 1.737 ;
      LAYER M5 ;
        RECT  24.882 1.057 25.002 29.723 ;
        RECT  18.978 1.057 19.098 29.723 ;
        RECT  13.074 1.057 13.194 29.723 ;
        RECT  7.17 1.057 7.29 29.723 ;
        RECT  1.266 1.057 1.386 29.723 ;
      LAYER M2 ;
        RECT  1.026 29.691 29.97 29.709 ;
        RECT  1.026 29.151 29.97 29.169 ;
        RECT  1.026 28.611 29.97 28.629 ;
        RECT  1.026 28.071 29.97 28.089 ;
        RECT  1.026 27.531 29.97 27.549 ;
        RECT  1.026 26.991 29.97 27.009 ;
        RECT  1.026 26.451 29.97 26.469 ;
        RECT  1.026 25.911 29.97 25.929 ;
        RECT  1.026 25.371 29.97 25.389 ;
        RECT  1.026 24.831 29.97 24.849 ;
        RECT  1.026 24.291 29.97 24.309 ;
        RECT  1.026 23.751 29.97 23.769 ;
        RECT  1.026 23.211 29.97 23.229 ;
        RECT  1.026 22.671 29.97 22.689 ;
        RECT  1.026 22.131 29.97 22.149 ;
        RECT  1.026 21.591 29.97 21.609 ;
        RECT  1.026 21.051 29.97 21.069 ;
        RECT  1.026 20.511 29.97 20.529 ;
        RECT  1.026 19.971 29.97 19.989 ;
        RECT  1.026 19.431 29.97 19.449 ;
        RECT  1.026 18.891 29.97 18.909 ;
        RECT  1.026 18.351 29.97 18.369 ;
        RECT  1.026 17.811 29.97 17.829 ;
        RECT  1.026 17.271 29.97 17.289 ;
        RECT  1.026 16.731 29.97 16.749 ;
        RECT  1.026 16.191 29.97 16.209 ;
        RECT  1.026 15.651 29.97 15.669 ;
        RECT  1.026 15.111 29.97 15.129 ;
        RECT  1.026 14.571 29.97 14.589 ;
        RECT  1.026 14.031 29.97 14.049 ;
        RECT  1.026 13.491 29.97 13.509 ;
        RECT  1.026 12.951 29.97 12.969 ;
        RECT  1.026 12.411 29.97 12.429 ;
        RECT  1.026 11.871 29.97 11.889 ;
        RECT  1.026 11.331 29.97 11.349 ;
        RECT  1.026 10.791 29.97 10.809 ;
        RECT  1.026 10.251 29.97 10.269 ;
        RECT  1.026 9.711 29.97 9.729 ;
        RECT  1.026 9.171 29.97 9.189 ;
        RECT  1.026 8.631 29.97 8.649 ;
        RECT  1.026 8.091 29.97 8.109 ;
        RECT  1.026 7.551 29.97 7.569 ;
        RECT  1.026 7.011 29.97 7.029 ;
        RECT  1.026 6.471 29.97 6.489 ;
        RECT  1.026 5.931 29.97 5.949 ;
        RECT  1.026 5.391 29.97 5.409 ;
        RECT  1.026 4.851 29.97 4.869 ;
        RECT  1.026 4.311 29.97 4.329 ;
        RECT  1.026 3.771 29.97 3.789 ;
        RECT  1.026 3.231 29.97 3.249 ;
        RECT  1.026 2.691 29.97 2.709 ;
        RECT  1.026 2.151 29.97 2.169 ;
        RECT  1.026 1.611 29.97 1.629 ;
        RECT  1.026 1.071 29.97 1.089 ;
      LAYER M1 ;
        RECT  1.026 29.691 29.97 29.709 ;
        RECT  1.026 29.151 29.97 29.169 ;
        RECT  1.026 28.611 29.97 28.629 ;
        RECT  1.026 28.071 29.97 28.089 ;
        RECT  1.026 27.531 29.97 27.549 ;
        RECT  1.026 26.991 29.97 27.009 ;
        RECT  1.026 26.451 29.97 26.469 ;
        RECT  1.026 25.911 29.97 25.929 ;
        RECT  1.026 25.371 29.97 25.389 ;
        RECT  1.026 24.831 29.97 24.849 ;
        RECT  1.026 24.291 29.97 24.309 ;
        RECT  1.026 23.751 29.97 23.769 ;
        RECT  1.026 23.211 29.97 23.229 ;
        RECT  1.026 22.671 29.97 22.689 ;
        RECT  1.026 22.131 29.97 22.149 ;
        RECT  1.026 21.591 29.97 21.609 ;
        RECT  1.026 21.051 29.97 21.069 ;
        RECT  1.026 20.511 29.97 20.529 ;
        RECT  1.026 19.971 29.97 19.989 ;
        RECT  1.026 19.431 29.97 19.449 ;
        RECT  1.026 18.891 29.97 18.909 ;
        RECT  1.026 18.351 29.97 18.369 ;
        RECT  1.026 17.811 29.97 17.829 ;
        RECT  1.026 17.271 29.97 17.289 ;
        RECT  1.026 16.731 29.97 16.749 ;
        RECT  1.026 16.191 29.97 16.209 ;
        RECT  1.026 15.651 29.97 15.669 ;
        RECT  1.026 15.111 29.97 15.129 ;
        RECT  1.026 14.571 29.97 14.589 ;
        RECT  1.026 14.031 29.97 14.049 ;
        RECT  1.026 13.491 29.97 13.509 ;
        RECT  1.026 12.951 29.97 12.969 ;
        RECT  1.026 12.411 29.97 12.429 ;
        RECT  1.026 11.871 29.97 11.889 ;
        RECT  1.026 11.331 29.97 11.349 ;
        RECT  1.026 10.791 29.97 10.809 ;
        RECT  1.026 10.251 29.97 10.269 ;
        RECT  1.026 9.711 29.97 9.729 ;
        RECT  1.026 9.171 29.97 9.189 ;
        RECT  1.026 8.631 29.97 8.649 ;
        RECT  1.026 8.091 29.97 8.109 ;
        RECT  1.026 7.551 29.97 7.569 ;
        RECT  1.026 7.011 29.97 7.029 ;
        RECT  1.026 6.471 29.97 6.489 ;
        RECT  1.026 5.931 29.97 5.949 ;
        RECT  1.026 5.391 29.97 5.409 ;
        RECT  1.026 4.851 29.97 4.869 ;
        RECT  1.026 4.311 29.97 4.329 ;
        RECT  1.026 3.771 29.97 3.789 ;
        RECT  1.026 3.231 29.97 3.249 ;
        RECT  1.026 2.691 29.97 2.709 ;
        RECT  1.026 2.151 29.97 2.169 ;
        RECT  1.026 1.611 29.97 1.629 ;
        RECT  1.026 1.071 29.97 1.089 ;
      VIA 24.942 25.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 19.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 13.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 7.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 1.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 25.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 19.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 13.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 7.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 1.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 25.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 19.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 13.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 7.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 1.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 25.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 19.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 13.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 7.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 1.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 25.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 19.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 13.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 7.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 1.593 CSRFile_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 29.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.683 24.987 29.717 ;
      VIA 24.942 29.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 29.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 29.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.143 24.987 29.177 ;
      VIA 24.942 29.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 29.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 28.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.603 24.987 28.637 ;
      VIA 24.942 28.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 28.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 28.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.063 24.987 28.097 ;
      VIA 24.942 28.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 28.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 27.54 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 27.523 24.987 27.557 ;
      VIA 24.942 27.54 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 27.54 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.983 24.987 27.017 ;
      VIA 24.942 27 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 27 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 26.46 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.443 24.987 26.477 ;
      VIA 24.942 26.46 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 26.46 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 25.92 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.903 24.987 25.937 ;
      VIA 24.942 25.92 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 25.92 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 25.38 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.363 24.987 25.397 ;
      VIA 24.942 25.38 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 25.38 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 24.84 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.823 24.987 24.857 ;
      VIA 24.942 24.84 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 24.84 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 24.3 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.283 24.987 24.317 ;
      VIA 24.942 24.3 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 24.3 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 23.76 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.743 24.987 23.777 ;
      VIA 24.942 23.76 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 23.76 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 23.22 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.203 24.987 23.237 ;
      VIA 24.942 23.22 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 23.22 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 22.68 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.663 24.987 22.697 ;
      VIA 24.942 22.68 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 22.68 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 22.14 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.123 24.987 22.157 ;
      VIA 24.942 22.14 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 22.14 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 21.6 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.583 24.987 21.617 ;
      VIA 24.942 21.6 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 21.6 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 21.06 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.043 24.987 21.077 ;
      VIA 24.942 21.06 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 21.06 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 20.52 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 20.503 24.987 20.537 ;
      VIA 24.942 20.52 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 20.52 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 19.98 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.963 24.987 19.997 ;
      VIA 24.942 19.98 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 19.98 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 19.44 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.423 24.987 19.457 ;
      VIA 24.942 19.44 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 19.44 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 18.9 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.883 24.987 18.917 ;
      VIA 24.942 18.9 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 18.9 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 18.36 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.343 24.987 18.377 ;
      VIA 24.942 18.36 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 18.36 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 17.82 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.803 24.987 17.837 ;
      VIA 24.942 17.82 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 17.82 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 17.28 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.263 24.987 17.297 ;
      VIA 24.942 17.28 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 17.28 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 16.74 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.723 24.987 16.757 ;
      VIA 24.942 16.74 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 16.74 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 16.2 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.183 24.987 16.217 ;
      VIA 24.942 16.2 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 16.2 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 15.66 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.643 24.987 15.677 ;
      VIA 24.942 15.66 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 15.66 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 15.12 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.103 24.987 15.137 ;
      VIA 24.942 15.12 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 15.12 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 14.58 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.563 24.987 14.597 ;
      VIA 24.942 14.58 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 14.58 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 14.04 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.023 24.987 14.057 ;
      VIA 24.942 14.04 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 14.04 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 13.5 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 13.483 24.987 13.517 ;
      VIA 24.942 13.5 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 13.5 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 12.96 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.943 24.987 12.977 ;
      VIA 24.942 12.96 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 12.96 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 12.42 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.403 24.987 12.437 ;
      VIA 24.942 12.42 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 12.42 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 11.88 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.863 24.987 11.897 ;
      VIA 24.942 11.88 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 11.88 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 11.34 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.323 24.987 11.357 ;
      VIA 24.942 11.34 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 11.34 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 10.8 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.783 24.987 10.817 ;
      VIA 24.942 10.8 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 10.8 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 10.26 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.243 24.987 10.277 ;
      VIA 24.942 10.26 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 10.26 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 9.72 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.703 24.987 9.737 ;
      VIA 24.942 9.72 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 9.72 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 9.18 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.163 24.987 9.197 ;
      VIA 24.942 9.18 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 9.18 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 8.64 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.623 24.987 8.657 ;
      VIA 24.942 8.64 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 8.64 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 8.1 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.083 24.987 8.117 ;
      VIA 24.942 8.1 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 8.1 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 7.56 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.543 24.987 7.577 ;
      VIA 24.942 7.56 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 7.56 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 7.02 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.003 24.987 7.037 ;
      VIA 24.942 7.02 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 7.02 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 6.48 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 6.463 24.987 6.497 ;
      VIA 24.942 6.48 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 6.48 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 5.94 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.923 24.987 5.957 ;
      VIA 24.942 5.94 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 5.94 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 5.4 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.383 24.987 5.417 ;
      VIA 24.942 5.4 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 5.4 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 4.86 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.843 24.987 4.877 ;
      VIA 24.942 4.86 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 4.86 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 4.32 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.303 24.987 4.337 ;
      VIA 24.942 4.32 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 4.32 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 3.78 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.763 24.987 3.797 ;
      VIA 24.942 3.78 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 3.78 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 3.24 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.223 24.987 3.257 ;
      VIA 24.942 3.24 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 3.24 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 2.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.683 24.987 2.717 ;
      VIA 24.942 2.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 2.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 2.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.143 24.987 2.177 ;
      VIA 24.942 2.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 2.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 1.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.603 24.987 1.637 ;
      VIA 24.942 1.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 1.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 24.942 1.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.063 24.987 1.097 ;
      VIA 24.942 1.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 24.942 1.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 29.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.683 19.083 29.717 ;
      VIA 19.038 29.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 29.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 29.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.143 19.083 29.177 ;
      VIA 19.038 29.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 29.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 28.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.603 19.083 28.637 ;
      VIA 19.038 28.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 28.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 28.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.063 19.083 28.097 ;
      VIA 19.038 28.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 28.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 27.54 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 27.523 19.083 27.557 ;
      VIA 19.038 27.54 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 27.54 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.983 19.083 27.017 ;
      VIA 19.038 27 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 27 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 26.46 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.443 19.083 26.477 ;
      VIA 19.038 26.46 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 26.46 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 25.92 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.903 19.083 25.937 ;
      VIA 19.038 25.92 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 25.92 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 25.38 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.363 19.083 25.397 ;
      VIA 19.038 25.38 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 25.38 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 24.84 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.823 19.083 24.857 ;
      VIA 19.038 24.84 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 24.84 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 24.3 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.283 19.083 24.317 ;
      VIA 19.038 24.3 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 24.3 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 23.76 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.743 19.083 23.777 ;
      VIA 19.038 23.76 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 23.76 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 23.22 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.203 19.083 23.237 ;
      VIA 19.038 23.22 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 23.22 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 22.68 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.663 19.083 22.697 ;
      VIA 19.038 22.68 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 22.68 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 22.14 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.123 19.083 22.157 ;
      VIA 19.038 22.14 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 22.14 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 21.6 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.583 19.083 21.617 ;
      VIA 19.038 21.6 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 21.6 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 21.06 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.043 19.083 21.077 ;
      VIA 19.038 21.06 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 21.06 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 20.52 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 20.503 19.083 20.537 ;
      VIA 19.038 20.52 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 20.52 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 19.98 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.963 19.083 19.997 ;
      VIA 19.038 19.98 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 19.98 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 19.44 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.423 19.083 19.457 ;
      VIA 19.038 19.44 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 19.44 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 18.9 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.883 19.083 18.917 ;
      VIA 19.038 18.9 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 18.9 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 18.36 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.343 19.083 18.377 ;
      VIA 19.038 18.36 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 18.36 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 17.82 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.803 19.083 17.837 ;
      VIA 19.038 17.82 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 17.82 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 17.28 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.263 19.083 17.297 ;
      VIA 19.038 17.28 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 17.28 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 16.74 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.723 19.083 16.757 ;
      VIA 19.038 16.74 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 16.74 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 16.2 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.183 19.083 16.217 ;
      VIA 19.038 16.2 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 16.2 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 15.66 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.643 19.083 15.677 ;
      VIA 19.038 15.66 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 15.66 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 15.12 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.103 19.083 15.137 ;
      VIA 19.038 15.12 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 15.12 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 14.58 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.563 19.083 14.597 ;
      VIA 19.038 14.58 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 14.58 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 14.04 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.023 19.083 14.057 ;
      VIA 19.038 14.04 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 14.04 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 13.5 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 13.483 19.083 13.517 ;
      VIA 19.038 13.5 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 13.5 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 12.96 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.943 19.083 12.977 ;
      VIA 19.038 12.96 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 12.96 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 12.42 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.403 19.083 12.437 ;
      VIA 19.038 12.42 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 12.42 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 11.88 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.863 19.083 11.897 ;
      VIA 19.038 11.88 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 11.88 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 11.34 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.323 19.083 11.357 ;
      VIA 19.038 11.34 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 11.34 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 10.8 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.783 19.083 10.817 ;
      VIA 19.038 10.8 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 10.8 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 10.26 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.243 19.083 10.277 ;
      VIA 19.038 10.26 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 10.26 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 9.72 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.703 19.083 9.737 ;
      VIA 19.038 9.72 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 9.72 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 9.18 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.163 19.083 9.197 ;
      VIA 19.038 9.18 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 9.18 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 8.64 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.623 19.083 8.657 ;
      VIA 19.038 8.64 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 8.64 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 8.1 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.083 19.083 8.117 ;
      VIA 19.038 8.1 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 8.1 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 7.56 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.543 19.083 7.577 ;
      VIA 19.038 7.56 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 7.56 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 7.02 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.003 19.083 7.037 ;
      VIA 19.038 7.02 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 7.02 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 6.48 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 6.463 19.083 6.497 ;
      VIA 19.038 6.48 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 6.48 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 5.94 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.923 19.083 5.957 ;
      VIA 19.038 5.94 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 5.94 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 5.4 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.383 19.083 5.417 ;
      VIA 19.038 5.4 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 5.4 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 4.86 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.843 19.083 4.877 ;
      VIA 19.038 4.86 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 4.86 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 4.32 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.303 19.083 4.337 ;
      VIA 19.038 4.32 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 4.32 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 3.78 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.763 19.083 3.797 ;
      VIA 19.038 3.78 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 3.78 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 3.24 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.223 19.083 3.257 ;
      VIA 19.038 3.24 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 3.24 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 2.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.683 19.083 2.717 ;
      VIA 19.038 2.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 2.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 2.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.143 19.083 2.177 ;
      VIA 19.038 2.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 2.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 1.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.603 19.083 1.637 ;
      VIA 19.038 1.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 1.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 19.038 1.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.063 19.083 1.097 ;
      VIA 19.038 1.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 19.038 1.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 29.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.683 13.179 29.717 ;
      VIA 13.134 29.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 29.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 29.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.143 13.179 29.177 ;
      VIA 13.134 29.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 29.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 28.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.603 13.179 28.637 ;
      VIA 13.134 28.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 28.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 28.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.063 13.179 28.097 ;
      VIA 13.134 28.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 28.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 27.54 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 27.523 13.179 27.557 ;
      VIA 13.134 27.54 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 27.54 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.983 13.179 27.017 ;
      VIA 13.134 27 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 27 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 26.46 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.443 13.179 26.477 ;
      VIA 13.134 26.46 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 26.46 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 25.92 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.903 13.179 25.937 ;
      VIA 13.134 25.92 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 25.92 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 25.38 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.363 13.179 25.397 ;
      VIA 13.134 25.38 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 25.38 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 24.84 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.823 13.179 24.857 ;
      VIA 13.134 24.84 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 24.84 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 24.3 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.283 13.179 24.317 ;
      VIA 13.134 24.3 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 24.3 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 23.76 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.743 13.179 23.777 ;
      VIA 13.134 23.76 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 23.76 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 23.22 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.203 13.179 23.237 ;
      VIA 13.134 23.22 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 23.22 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 22.68 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.663 13.179 22.697 ;
      VIA 13.134 22.68 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 22.68 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 22.14 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.123 13.179 22.157 ;
      VIA 13.134 22.14 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 22.14 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 21.6 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.583 13.179 21.617 ;
      VIA 13.134 21.6 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 21.6 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 21.06 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.043 13.179 21.077 ;
      VIA 13.134 21.06 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 21.06 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 20.52 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 20.503 13.179 20.537 ;
      VIA 13.134 20.52 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 20.52 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 19.98 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.963 13.179 19.997 ;
      VIA 13.134 19.98 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 19.98 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 19.44 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.423 13.179 19.457 ;
      VIA 13.134 19.44 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 19.44 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 18.9 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.883 13.179 18.917 ;
      VIA 13.134 18.9 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 18.9 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 18.36 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.343 13.179 18.377 ;
      VIA 13.134 18.36 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 18.36 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 17.82 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.803 13.179 17.837 ;
      VIA 13.134 17.82 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 17.82 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 17.28 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.263 13.179 17.297 ;
      VIA 13.134 17.28 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 17.28 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 16.74 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.723 13.179 16.757 ;
      VIA 13.134 16.74 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 16.74 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 16.2 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.183 13.179 16.217 ;
      VIA 13.134 16.2 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 16.2 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 15.66 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.643 13.179 15.677 ;
      VIA 13.134 15.66 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 15.66 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 15.12 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.103 13.179 15.137 ;
      VIA 13.134 15.12 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 15.12 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 14.58 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.563 13.179 14.597 ;
      VIA 13.134 14.58 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 14.58 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 14.04 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.023 13.179 14.057 ;
      VIA 13.134 14.04 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 14.04 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 13.5 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 13.483 13.179 13.517 ;
      VIA 13.134 13.5 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 13.5 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 12.96 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.943 13.179 12.977 ;
      VIA 13.134 12.96 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 12.96 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 12.42 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.403 13.179 12.437 ;
      VIA 13.134 12.42 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 12.42 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 11.88 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.863 13.179 11.897 ;
      VIA 13.134 11.88 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 11.88 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 11.34 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.323 13.179 11.357 ;
      VIA 13.134 11.34 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 11.34 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 10.8 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.783 13.179 10.817 ;
      VIA 13.134 10.8 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 10.8 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 10.26 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.243 13.179 10.277 ;
      VIA 13.134 10.26 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 10.26 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 9.72 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.703 13.179 9.737 ;
      VIA 13.134 9.72 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 9.72 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 9.18 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.163 13.179 9.197 ;
      VIA 13.134 9.18 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 9.18 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 8.64 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.623 13.179 8.657 ;
      VIA 13.134 8.64 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 8.64 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 8.1 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.083 13.179 8.117 ;
      VIA 13.134 8.1 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 8.1 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 7.56 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.543 13.179 7.577 ;
      VIA 13.134 7.56 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 7.56 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 7.02 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.003 13.179 7.037 ;
      VIA 13.134 7.02 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 7.02 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 6.48 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 6.463 13.179 6.497 ;
      VIA 13.134 6.48 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 6.48 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 5.94 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.923 13.179 5.957 ;
      VIA 13.134 5.94 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 5.94 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 5.4 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.383 13.179 5.417 ;
      VIA 13.134 5.4 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 5.4 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 4.86 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.843 13.179 4.877 ;
      VIA 13.134 4.86 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 4.86 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 4.32 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.303 13.179 4.337 ;
      VIA 13.134 4.32 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 4.32 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 3.78 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.763 13.179 3.797 ;
      VIA 13.134 3.78 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 3.78 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 3.24 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.223 13.179 3.257 ;
      VIA 13.134 3.24 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 3.24 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 2.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.683 13.179 2.717 ;
      VIA 13.134 2.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 2.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 2.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.143 13.179 2.177 ;
      VIA 13.134 2.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 2.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 1.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.603 13.179 1.637 ;
      VIA 13.134 1.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 1.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 13.134 1.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.063 13.179 1.097 ;
      VIA 13.134 1.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 13.134 1.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 29.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.683 7.275 29.717 ;
      VIA 7.23 29.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 29.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 29.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.143 7.275 29.177 ;
      VIA 7.23 29.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 29.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 28.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.603 7.275 28.637 ;
      VIA 7.23 28.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 28.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 28.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.063 7.275 28.097 ;
      VIA 7.23 28.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 28.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 27.54 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 27.523 7.275 27.557 ;
      VIA 7.23 27.54 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 27.54 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.983 7.275 27.017 ;
      VIA 7.23 27 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 27 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 26.46 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.443 7.275 26.477 ;
      VIA 7.23 26.46 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 26.46 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 25.92 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.903 7.275 25.937 ;
      VIA 7.23 25.92 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 25.92 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 25.38 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.363 7.275 25.397 ;
      VIA 7.23 25.38 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 25.38 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 24.84 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.823 7.275 24.857 ;
      VIA 7.23 24.84 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 24.84 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 24.3 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.283 7.275 24.317 ;
      VIA 7.23 24.3 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 24.3 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 23.76 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.743 7.275 23.777 ;
      VIA 7.23 23.76 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 23.76 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 23.22 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.203 7.275 23.237 ;
      VIA 7.23 23.22 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 23.22 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 22.68 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.663 7.275 22.697 ;
      VIA 7.23 22.68 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 22.68 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 22.14 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.123 7.275 22.157 ;
      VIA 7.23 22.14 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 22.14 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 21.6 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.583 7.275 21.617 ;
      VIA 7.23 21.6 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 21.6 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 21.06 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.043 7.275 21.077 ;
      VIA 7.23 21.06 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 21.06 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 20.52 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 20.503 7.275 20.537 ;
      VIA 7.23 20.52 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 20.52 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 19.98 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.963 7.275 19.997 ;
      VIA 7.23 19.98 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 19.98 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 19.44 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.423 7.275 19.457 ;
      VIA 7.23 19.44 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 19.44 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 18.9 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.883 7.275 18.917 ;
      VIA 7.23 18.9 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 18.9 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 18.36 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.343 7.275 18.377 ;
      VIA 7.23 18.36 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 18.36 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 17.82 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.803 7.275 17.837 ;
      VIA 7.23 17.82 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 17.82 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 17.28 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.263 7.275 17.297 ;
      VIA 7.23 17.28 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 17.28 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 16.74 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.723 7.275 16.757 ;
      VIA 7.23 16.74 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 16.74 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 16.2 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.183 7.275 16.217 ;
      VIA 7.23 16.2 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 16.2 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 15.66 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.643 7.275 15.677 ;
      VIA 7.23 15.66 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 15.66 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 15.12 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.103 7.275 15.137 ;
      VIA 7.23 15.12 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 15.12 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 14.58 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.563 7.275 14.597 ;
      VIA 7.23 14.58 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 14.58 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 14.04 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.023 7.275 14.057 ;
      VIA 7.23 14.04 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 14.04 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 13.5 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 13.483 7.275 13.517 ;
      VIA 7.23 13.5 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 13.5 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 12.96 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.943 7.275 12.977 ;
      VIA 7.23 12.96 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 12.96 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 12.42 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.403 7.275 12.437 ;
      VIA 7.23 12.42 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 12.42 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 11.88 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.863 7.275 11.897 ;
      VIA 7.23 11.88 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 11.88 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 11.34 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.323 7.275 11.357 ;
      VIA 7.23 11.34 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 11.34 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 10.8 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.783 7.275 10.817 ;
      VIA 7.23 10.8 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 10.8 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 10.26 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.243 7.275 10.277 ;
      VIA 7.23 10.26 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 10.26 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 9.72 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.703 7.275 9.737 ;
      VIA 7.23 9.72 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 9.72 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 9.18 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.163 7.275 9.197 ;
      VIA 7.23 9.18 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 9.18 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 8.64 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.623 7.275 8.657 ;
      VIA 7.23 8.64 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 8.64 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 8.1 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.083 7.275 8.117 ;
      VIA 7.23 8.1 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 8.1 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 7.56 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.543 7.275 7.577 ;
      VIA 7.23 7.56 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 7.56 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 7.02 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.003 7.275 7.037 ;
      VIA 7.23 7.02 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 7.02 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 6.48 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 6.463 7.275 6.497 ;
      VIA 7.23 6.48 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 6.48 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 5.94 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.923 7.275 5.957 ;
      VIA 7.23 5.94 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 5.94 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 5.4 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.383 7.275 5.417 ;
      VIA 7.23 5.4 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 5.4 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 4.86 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.843 7.275 4.877 ;
      VIA 7.23 4.86 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 4.86 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 4.32 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.303 7.275 4.337 ;
      VIA 7.23 4.32 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 4.32 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 3.78 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.763 7.275 3.797 ;
      VIA 7.23 3.78 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 3.78 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 3.24 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.223 7.275 3.257 ;
      VIA 7.23 3.24 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 3.24 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 2.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.683 7.275 2.717 ;
      VIA 7.23 2.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 2.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 2.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.143 7.275 2.177 ;
      VIA 7.23 2.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 2.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 1.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.603 7.275 1.637 ;
      VIA 7.23 1.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 1.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 7.23 1.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.063 7.275 1.097 ;
      VIA 7.23 1.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 7.23 1.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 29.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.683 1.371 29.717 ;
      VIA 1.326 29.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 29.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 29.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.143 1.371 29.177 ;
      VIA 1.326 29.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 29.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 28.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.603 1.371 28.637 ;
      VIA 1.326 28.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 28.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 28.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.063 1.371 28.097 ;
      VIA 1.326 28.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 28.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 27.54 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 27.523 1.371 27.557 ;
      VIA 1.326 27.54 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 27.54 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 27 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.983 1.371 27.017 ;
      VIA 1.326 27 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 27 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 26.46 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.443 1.371 26.477 ;
      VIA 1.326 26.46 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 26.46 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 25.92 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.903 1.371 25.937 ;
      VIA 1.326 25.92 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 25.92 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 25.38 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.363 1.371 25.397 ;
      VIA 1.326 25.38 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 25.38 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 24.84 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.823 1.371 24.857 ;
      VIA 1.326 24.84 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 24.84 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 24.3 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.283 1.371 24.317 ;
      VIA 1.326 24.3 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 24.3 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 23.76 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.743 1.371 23.777 ;
      VIA 1.326 23.76 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 23.76 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 23.22 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.203 1.371 23.237 ;
      VIA 1.326 23.22 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 23.22 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 22.68 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.663 1.371 22.697 ;
      VIA 1.326 22.68 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 22.68 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 22.14 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.123 1.371 22.157 ;
      VIA 1.326 22.14 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 22.14 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 21.6 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.583 1.371 21.617 ;
      VIA 1.326 21.6 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 21.6 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 21.06 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.043 1.371 21.077 ;
      VIA 1.326 21.06 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 21.06 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 20.52 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 20.503 1.371 20.537 ;
      VIA 1.326 20.52 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 20.52 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 19.98 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.963 1.371 19.997 ;
      VIA 1.326 19.98 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 19.98 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 19.44 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.423 1.371 19.457 ;
      VIA 1.326 19.44 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 19.44 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 18.9 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.883 1.371 18.917 ;
      VIA 1.326 18.9 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 18.9 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 18.36 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.343 1.371 18.377 ;
      VIA 1.326 18.36 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 18.36 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 17.82 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.803 1.371 17.837 ;
      VIA 1.326 17.82 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 17.82 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 17.28 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.263 1.371 17.297 ;
      VIA 1.326 17.28 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 17.28 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 16.74 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.723 1.371 16.757 ;
      VIA 1.326 16.74 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 16.74 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 16.2 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.183 1.371 16.217 ;
      VIA 1.326 16.2 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 16.2 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 15.66 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.643 1.371 15.677 ;
      VIA 1.326 15.66 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 15.66 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 15.12 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.103 1.371 15.137 ;
      VIA 1.326 15.12 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 15.12 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 14.58 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.563 1.371 14.597 ;
      VIA 1.326 14.58 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 14.58 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 14.04 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.023 1.371 14.057 ;
      VIA 1.326 14.04 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 14.04 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 13.5 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 13.483 1.371 13.517 ;
      VIA 1.326 13.5 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 13.5 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 12.96 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.943 1.371 12.977 ;
      VIA 1.326 12.96 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 12.96 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 12.42 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.403 1.371 12.437 ;
      VIA 1.326 12.42 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 12.42 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 11.88 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.863 1.371 11.897 ;
      VIA 1.326 11.88 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 11.88 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 11.34 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.323 1.371 11.357 ;
      VIA 1.326 11.34 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 11.34 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 10.8 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.783 1.371 10.817 ;
      VIA 1.326 10.8 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 10.8 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 10.26 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.243 1.371 10.277 ;
      VIA 1.326 10.26 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 10.26 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 9.72 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.703 1.371 9.737 ;
      VIA 1.326 9.72 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 9.72 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 9.18 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.163 1.371 9.197 ;
      VIA 1.326 9.18 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 9.18 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 8.64 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.623 1.371 8.657 ;
      VIA 1.326 8.64 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 8.64 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 8.1 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.083 1.371 8.117 ;
      VIA 1.326 8.1 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 8.1 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 7.56 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.543 1.371 7.577 ;
      VIA 1.326 7.56 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 7.56 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 7.02 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.003 1.371 7.037 ;
      VIA 1.326 7.02 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 7.02 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 6.48 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 6.463 1.371 6.497 ;
      VIA 1.326 6.48 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 6.48 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 5.94 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.923 1.371 5.957 ;
      VIA 1.326 5.94 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 5.94 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 5.4 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.383 1.371 5.417 ;
      VIA 1.326 5.4 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 5.4 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 4.86 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 CSRFile_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 CSRFile_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 CSRFile_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 CSRFile_VIA23_1_3_36_36 ;
      VIA 15.498 29.7 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 29.16 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 28.62 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 28.08 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 27.54 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 27 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 26.46 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 25.92 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 25.38 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 24.84 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 24.3 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 23.76 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 23.22 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 22.68 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 22.14 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 21.6 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 21.06 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 20.52 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 19.98 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 19.44 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 18.9 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 18.36 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 17.82 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 17.28 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 16.74 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 16.2 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 15.66 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 15.12 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 14.58 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 14.04 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 13.5 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 12.96 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 12.42 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 11.88 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 11.34 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 10.8 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 10.26 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 9.72 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 9.18 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 8.64 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 8.1 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 7.56 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 7.02 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 6.48 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 5.94 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 5.4 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 4.86 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 4.32 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 3.78 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 3.24 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 2.7 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 2.16 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 1.62 CSRFile_via1_2_28944_18_1_804_36_36 ;
      VIA 15.498 1.08 CSRFile_via1_2_28944_18_1_804_36_36 ;
    END
  END VSS
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 3.648 31.005 3.672 ;
    END
  END clock
  PIN io_cause[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.176 0 10.2 0.084 ;
    END
  END io_cause[0]
  PIN io_cause[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.288 0 12.312 0.084 ;
    END
  END io_cause[10]
  PIN io_cause[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.328 0 11.352 0.084 ;
    END
  END io_cause[11]
  PIN io_cause[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.464 0.084 10.488 ;
    END
  END io_cause[12]
  PIN io_cause[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.088 0.084 17.112 ;
    END
  END io_cause[13]
  PIN io_cause[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.528 0.084 18.552 ;
    END
  END io_cause[14]
  PIN io_cause[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.704 0.084 16.728 ;
    END
  END io_cause[15]
  PIN io_cause[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.776 0.084 19.8 ;
    END
  END io_cause[16]
  PIN io_cause[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.64 30.921 8.664 31.005 ;
    END
  END io_cause[17]
  PIN io_cause[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.752 0.084 22.776 ;
    END
  END io_cause[18]
  PIN io_cause[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.272 30.921 10.296 31.005 ;
    END
  END io_cause[19]
  PIN io_cause[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.968 0 7.992 0.084 ;
    END
  END io_cause[1]
  PIN io_cause[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.16 30.921 8.184 31.005 ;
    END
  END io_cause[20]
  PIN io_cause[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.464 30.921 10.488 31.005 ;
    END
  END io_cause[21]
  PIN io_cause[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.944 30.921 10.968 31.005 ;
    END
  END io_cause[22]
  PIN io_cause[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.68 30.921 7.704 31.005 ;
    END
  END io_cause[23]
  PIN io_cause[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.512 0.084 16.536 ;
    END
  END io_cause[24]
  PIN io_cause[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.872 0.084 19.896 ;
    END
  END io_cause[25]
  PIN io_cause[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.528 30.921 6.552 31.005 ;
    END
  END io_cause[26]
  PIN io_cause[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.024 0.084 21.048 ;
    END
  END io_cause[27]
  PIN io_cause[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.888 0.084 21.912 ;
    END
  END io_cause[28]
  PIN io_cause[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.472 0.084 17.496 ;
    END
  END io_cause[29]
  PIN io_cause[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 6.432 0.084 6.456 ;
    END
  END io_cause[2]
  PIN io_cause[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.376 0.084 17.4 ;
    END
  END io_cause[30]
  PIN io_cause[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.584 0.084 7.608 ;
    END
  END io_cause[31]
  PIN io_cause[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.488 0.084 7.512 ;
    END
  END io_cause[3]
  PIN io_cause[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 6.912 0.084 6.936 ;
    END
  END io_cause[4]
  PIN io_cause[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.832 0.084 8.856 ;
    END
  END io_cause[5]
  PIN io_cause[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.216 0.084 9.24 ;
    END
  END io_cause[6]
  PIN io_cause[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.256 0.084 8.28 ;
    END
  END io_cause[7]
  PIN io_cause[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.552 0.084 15.576 ;
    END
  END io_cause[8]
  PIN io_cause[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.304 0.084 14.328 ;
    END
  END io_cause[9]
  PIN io_eret
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.464 0 10.488 0.084 ;
    END
  END io_eret
  PIN io_evec[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.712 0 23.736 0.084 ;
    END
  END io_evec[0]
  PIN io_evec[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.608 0.084 16.632 ;
    END
  END io_evec[10]
  PIN io_evec[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.272 0 10.296 0.084 ;
    END
  END io_evec[11]
  PIN io_evec[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.56 0.084 10.584 ;
    END
  END io_evec[12]
  PIN io_evec[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.36 0.084 15.384 ;
    END
  END io_evec[13]
  PIN io_evec[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.624 0.084 18.648 ;
    END
  END io_evec[14]
  PIN io_evec[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.648 0.084 15.672 ;
    END
  END io_evec[15]
  PIN io_evec[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.392 0.084 19.416 ;
    END
  END io_evec[16]
  PIN io_evec[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.56 30.921 10.584 31.005 ;
    END
  END io_evec[17]
  PIN io_evec[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  5.76 30.921 5.784 31.005 ;
    END
  END io_evec[18]
  PIN io_evec[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.368 30.921 10.392 31.005 ;
    END
  END io_evec[19]
  PIN io_evec[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.616 0 23.64 0.084 ;
    END
  END io_evec[1]
  PIN io_evec[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.984 0.084 22.008 ;
    END
  END io_evec[20]
  PIN io_evec[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.112 30.921 14.136 31.005 ;
    END
  END io_evec[21]
  PIN io_evec[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.016 30.921 14.04 31.005 ;
    END
  END io_evec[22]
  PIN io_evec[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.544 30.921 8.568 31.005 ;
    END
  END io_evec[23]
  PIN io_evec[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.264 0.084 15.288 ;
    END
  END io_evec[24]
  PIN io_evec[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.16 0.084 20.184 ;
    END
  END io_evec[25]
  PIN io_evec[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.72 30.921 6.744 31.005 ;
    END
  END io_evec[26]
  PIN io_evec[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.64 0.084 20.664 ;
    END
  END io_evec[27]
  PIN io_evec[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.928 0.084 20.952 ;
    END
  END io_evec[28]
  PIN io_evec[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.184 0.084 17.208 ;
    END
  END io_evec[29]
  PIN io_evec[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.104 0.084 7.128 ;
    END
  END io_evec[2]
  PIN io_evec[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.816 0.084 18.84 ;
    END
  END io_evec[30]
  PIN io_evec[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.752 0 10.776 0.084 ;
    END
  END io_evec[31]
  PIN io_evec[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.832 0 8.856 0.084 ;
    END
  END io_evec[3]
  PIN io_evec[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.296 0.084 7.32 ;
    END
  END io_evec[4]
  PIN io_evec[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.392 0.084 7.416 ;
    END
  END io_evec[5]
  PIN io_evec[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.2 0.084 7.224 ;
    END
  END io_evec[6]
  PIN io_evec[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.152 0 13.176 0.084 ;
    END
  END io_evec[7]
  PIN io_evec[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.096 0 12.12 0.084 ;
    END
  END io_evec[8]
  PIN io_evec[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.536 0.084 13.56 ;
    END
  END io_evec[9]
  PIN io_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.112 0 14.136 0.084 ;
    END
  END io_exception
  PIN io_hartid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.128 0 16.152 0.084 ;
    END
  END io_hartid
  PIN io_interrupt
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.032 0 16.056 0.084 ;
    END
  END io_interrupt
  PIN io_interrupt_cause[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.208 0 14.232 0.084 ;
    END
  END io_interrupt_cause[0]
  PIN io_interrupt_cause[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.944 0 22.968 0.084 ;
    END
  END io_interrupt_cause[10]
  PIN io_interrupt_cause[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.272 0 22.296 0.084 ;
    END
  END io_interrupt_cause[11]
  PIN io_interrupt_cause[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.52 0 23.544 0.084 ;
    END
  END io_interrupt_cause[12]
  PIN io_interrupt_cause[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.504 0 21.528 0.084 ;
    END
  END io_interrupt_cause[13]
  PIN io_interrupt_cause[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.368 0 22.392 0.084 ;
    END
  END io_interrupt_cause[14]
  PIN io_interrupt_cause[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.888 0 21.912 0.084 ;
    END
  END io_interrupt_cause[15]
  PIN io_interrupt_cause[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.232 0 23.256 0.084 ;
    END
  END io_interrupt_cause[16]
  PIN io_interrupt_cause[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 0 21.72 0.084 ;
    END
  END io_interrupt_cause[17]
  PIN io_interrupt_cause[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.216 0 21.24 0.084 ;
    END
  END io_interrupt_cause[18]
  PIN io_interrupt_cause[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.408 0 21.432 0.084 ;
    END
  END io_interrupt_cause[19]
  PIN io_interrupt_cause[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.4 0 14.424 0.084 ;
    END
  END io_interrupt_cause[1]
  PIN io_interrupt_cause[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.464 0 22.488 0.084 ;
    END
  END io_interrupt_cause[20]
  PIN io_interrupt_cause[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.792 0 21.816 0.084 ;
    END
  END io_interrupt_cause[21]
  PIN io_interrupt_cause[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.848 0 22.872 0.084 ;
    END
  END io_interrupt_cause[22]
  PIN io_interrupt_cause[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.56 0 22.584 0.084 ;
    END
  END io_interrupt_cause[23]
  PIN io_interrupt_cause[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.12 0 21.144 0.084 ;
    END
  END io_interrupt_cause[24]
  PIN io_interrupt_cause[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.312 0 21.336 0.084 ;
    END
  END io_interrupt_cause[25]
  PIN io_interrupt_cause[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.024 0 21.048 0.084 ;
    END
  END io_interrupt_cause[26]
  PIN io_interrupt_cause[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.424 0 23.448 0.084 ;
    END
  END io_interrupt_cause[27]
  PIN io_interrupt_cause[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.752 0 22.776 0.084 ;
    END
  END io_interrupt_cause[28]
  PIN io_interrupt_cause[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.08 0 22.104 0.084 ;
    END
  END io_interrupt_cause[29]
  PIN io_interrupt_cause[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.016 0 14.04 0.084 ;
    END
  END io_interrupt_cause[2]
  PIN io_interrupt_cause[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.928 0 20.952 0.084 ;
    END
  END io_interrupt_cause[30]
  PIN io_interrupt_cause[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.728 30.921 1.752 31.005 ;
    END
  END io_interrupt_cause[31]
  PIN io_interrupt_cause[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.92 0 13.944 0.084 ;
    END
  END io_interrupt_cause[3]
  PIN io_interrupt_cause[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.136 0 23.16 0.084 ;
    END
  END io_interrupt_cause[4]
  PIN io_interrupt_cause[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.656 0 22.68 0.084 ;
    END
  END io_interrupt_cause[5]
  PIN io_interrupt_cause[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.328 0 23.352 0.084 ;
    END
  END io_interrupt_cause[6]
  PIN io_interrupt_cause[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.6 0 21.624 0.084 ;
    END
  END io_interrupt_cause[7]
  PIN io_interrupt_cause[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.176 0 22.2 0.084 ;
    END
  END io_interrupt_cause[8]
  PIN io_interrupt_cause[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.04 0 23.064 0.084 ;
    END
  END io_interrupt_cause[9]
  PIN io_interrupts_debug
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.248 0 13.272 0.084 ;
    END
  END io_interrupts_debug
  PIN io_interrupts_meip
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.672 0 12.696 0.084 ;
    END
  END io_interrupts_meip
  PIN io_interrupts_msip
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.344 0 13.368 0.084 ;
    END
  END io_interrupts_msip
  PIN io_interrupts_mtip
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.056 0 13.08 0.084 ;
    END
  END io_interrupts_mtip
  PIN io_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.672 0 0.696 0.084 ;
    END
  END io_pc[0]
  PIN io_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.128 0.084 16.152 ;
    END
  END io_pc[10]
  PIN io_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.312 0 9.336 0.084 ;
    END
  END io_pc[11]
  PIN io_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.752 0.084 10.776 ;
    END
  END io_pc[12]
  PIN io_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.936 0.084 15.96 ;
    END
  END io_pc[13]
  PIN io_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.048 0.084 18.072 ;
    END
  END io_pc[14]
  PIN io_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.576 0 12.6 0.084 ;
    END
  END io_pc[15]
  PIN io_pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.336 0.084 18.36 ;
    END
  END io_pc[16]
  PIN io_pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.216 30.921 9.24 31.005 ;
    END
  END io_pc[17]
  PIN io_pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.616 0.084 23.64 ;
    END
  END io_pc[18]
  PIN io_pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.656 30.921 10.68 31.005 ;
    END
  END io_pc[19]
  PIN io_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.768 0 0.792 0.084 ;
    END
  END io_pc[1]
  PIN io_pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.464 0.084 22.488 ;
    END
  END io_pc[20]
  PIN io_pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.848 30.921 10.872 31.005 ;
    END
  END io_pc[21]
  PIN io_pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.04 0.084 23.064 ;
    END
  END io_pc[22]
  PIN io_pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.488 30.921 7.512 31.005 ;
    END
  END io_pc[23]
  PIN io_pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.4 0.084 14.424 ;
    END
  END io_pc[24]
  PIN io_pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.312 0.084 21.336 ;
    END
  END io_pc[25]
  PIN io_pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  5.568 30.921 5.592 31.005 ;
    END
  END io_pc[26]
  PIN io_pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.544 0.084 20.568 ;
    END
  END io_pc[27]
  PIN io_pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.448 0.084 20.472 ;
    END
  END io_pc[28]
  PIN io_pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.992 0.084 17.016 ;
    END
  END io_pc[29]
  PIN io_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.448 0.084 8.472 ;
    END
  END io_pc[2]
  PIN io_pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.104 0.084 19.128 ;
    END
  END io_pc[30]
  PIN io_pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.024 0 9.048 0.084 ;
    END
  END io_pc[31]
  PIN io_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.928 0.084 8.952 ;
    END
  END io_pc[3]
  PIN io_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.544 0.084 8.568 ;
    END
  END io_pc[4]
  PIN io_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.656 0.084 10.68 ;
    END
  END io_pc[5]
  PIN io_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.176 0.084 10.2 ;
    END
  END io_pc[6]
  PIN io_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.616 0 11.64 0.084 ;
    END
  END io_pc[7]
  PIN io_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.656 0 10.68 0.084 ;
    END
  END io_pc[8]
  PIN io_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.728 0.084 13.752 ;
    END
  END io_pc[9]
  PIN io_retire
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 0 22.008 0.084 ;
    END
  END io_retire
  PIN io_rw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.864 0 12.888 0.084 ;
    END
  END io_rw_addr[0]
  PIN io_rw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.936 0 15.96 0.084 ;
    END
  END io_rw_addr[10]
  PIN io_rw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.648 0 15.672 0.084 ;
    END
  END io_rw_addr[11]
  PIN io_rw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.768 0 12.792 0.084 ;
    END
  END io_rw_addr[1]
  PIN io_rw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.304 0 14.328 0.084 ;
    END
  END io_rw_addr[2]
  PIN io_rw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.536 0 13.56 0.084 ;
    END
  END io_rw_addr[3]
  PIN io_rw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.84 0 15.864 0.084 ;
    END
  END io_rw_addr[4]
  PIN io_rw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.552 0 15.576 0.084 ;
    END
  END io_rw_addr[5]
  PIN io_rw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.44 0 13.464 0.084 ;
    END
  END io_rw_addr[6]
  PIN io_rw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.744 0 15.768 0.084 ;
    END
  END io_rw_addr[7]
  PIN io_rw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.456 0 15.48 0.084 ;
    END
  END io_rw_addr[8]
  PIN io_rw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.496 0 14.52 0.084 ;
    END
  END io_rw_addr[9]
  PIN io_rw_cmd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.224 0 16.248 0.084 ;
    END
  END io_rw_cmd[0]
  PIN io_rw_cmd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.32 0 16.344 0.084 ;
    END
  END io_rw_cmd[1]
  PIN io_rw_cmd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.416 0 16.44 0.084 ;
    END
  END io_rw_cmd[2]
  PIN io_rw_rdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.608 0 16.632 0.084 ;
    END
  END io_rw_rdata[0]
  PIN io_rw_rdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.976 0 15 0.084 ;
    END
  END io_rw_rdata[10]
  PIN io_rw_rdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.824 0 13.848 0.084 ;
    END
  END io_rw_rdata[11]
  PIN io_rw_rdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.88 0 14.904 0.084 ;
    END
  END io_rw_rdata[12]
  PIN io_rw_rdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.84 0.084 15.864 ;
    END
  END io_rw_rdata[13]
  PIN io_rw_rdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.432 30.921 18.456 31.005 ;
    END
  END io_rw_rdata[14]
  PIN io_rw_rdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.456 0.084 15.48 ;
    END
  END io_rw_rdata[15]
  PIN io_rw_rdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.72 0.084 18.744 ;
    END
  END io_rw_rdata[16]
  PIN io_rw_rdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.008 30.921 19.032 31.005 ;
    END
  END io_rw_rdata[17]
  PIN io_rw_rdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.592 30.921 14.616 31.005 ;
    END
  END io_rw_rdata[18]
  PIN io_rw_rdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.456 30.921 15.48 31.005 ;
    END
  END io_rw_rdata[19]
  PIN io_rw_rdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.832 0 20.856 0.084 ;
    END
  END io_rw_rdata[1]
  PIN io_rw_rdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.168 30.921 15.192 31.005 ;
    END
  END io_rw_rdata[20]
  PIN io_rw_rdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.36 30.921 15.384 31.005 ;
    END
  END io_rw_rdata[21]
  PIN io_rw_rdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.784 30.921 14.808 31.005 ;
    END
  END io_rw_rdata[22]
  PIN io_rw_rdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.128 30.921 16.152 31.005 ;
    END
  END io_rw_rdata[23]
  PIN io_rw_rdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.8 0.084 16.824 ;
    END
  END io_rw_rdata[24]
  PIN io_rw_rdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.736 0.084 20.76 ;
    END
  END io_rw_rdata[25]
  PIN io_rw_rdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.744 30.921 15.768 31.005 ;
    END
  END io_rw_rdata[26]
  PIN io_rw_rdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.256 0.084 20.28 ;
    END
  END io_rw_rdata[27]
  PIN io_rw_rdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.912 30.921 18.936 31.005 ;
    END
  END io_rw_rdata[28]
  PIN io_rw_rdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.568 0.084 17.592 ;
    END
  END io_rw_rdata[29]
  PIN io_rw_rdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.16 0 20.184 0.084 ;
    END
  END io_rw_rdata[2]
  PIN io_rw_rdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.432 0.084 18.456 ;
    END
  END io_rw_rdata[30]
  PIN io_rw_rdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 12.288 31.005 12.312 ;
    END
  END io_rw_rdata[31]
  PIN io_rw_rdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.992 0 17.016 0.084 ;
    END
  END io_rw_rdata[3]
  PIN io_rw_rdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.968 0 19.992 0.084 ;
    END
  END io_rw_rdata[4]
  PIN io_rw_rdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.192 0 12.216 0.084 ;
    END
  END io_rw_rdata[5]
  PIN io_rw_rdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 9.216 31.005 9.24 ;
    END
  END io_rw_rdata[6]
  PIN io_rw_rdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.28 0 17.304 0.084 ;
    END
  END io_rw_rdata[7]
  PIN io_rw_rdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.264 0 15.288 0.084 ;
    END
  END io_rw_rdata[8]
  PIN io_rw_rdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.168 0 15.192 0.084 ;
    END
  END io_rw_rdata[9]
  PIN io_rw_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.512 0 16.536 0.084 ;
    END
  END io_rw_wdata[0]
  PIN io_rw_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.688 0 14.712 0.084 ;
    END
  END io_rw_wdata[10]
  PIN io_rw_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.632 0 13.656 0.084 ;
    END
  END io_rw_wdata[11]
  PIN io_rw_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.592 0 14.616 0.084 ;
    END
  END io_rw_wdata[12]
  PIN io_rw_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.36 0 15.384 0.084 ;
    END
  END io_rw_wdata[13]
  PIN io_rw_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.336 30.921 18.36 31.005 ;
    END
  END io_rw_wdata[14]
  PIN io_rw_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.744 0.084 15.768 ;
    END
  END io_rw_wdata[15]
  PIN io_rw_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.008 0.084 19.032 ;
    END
  END io_rw_wdata[16]
  PIN io_rw_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.816 30.921 18.84 31.005 ;
    END
  END io_rw_wdata[17]
  PIN io_rw_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.976 30.921 15 31.005 ;
    END
  END io_rw_wdata[18]
  PIN io_rw_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.264 30.921 15.288 31.005 ;
    END
  END io_rw_wdata[19]
  PIN io_rw_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.448 0 20.472 0.084 ;
    END
  END io_rw_wdata[1]
  PIN io_rw_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.88 30.921 14.904 31.005 ;
    END
  END io_rw_wdata[20]
  PIN io_rw_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.072 30.921 15.096 31.005 ;
    END
  END io_rw_wdata[21]
  PIN io_rw_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.688 30.921 14.712 31.005 ;
    END
  END io_rw_wdata[22]
  PIN io_rw_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.84 30.921 15.864 31.005 ;
    END
  END io_rw_wdata[23]
  PIN io_rw_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.896 0.084 16.92 ;
    END
  END io_rw_wdata[24]
  PIN io_rw_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.832 0.084 20.856 ;
    END
  END io_rw_wdata[25]
  PIN io_rw_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.552 30.921 15.576 31.005 ;
    END
  END io_rw_wdata[26]
  PIN io_rw_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.064 0.084 20.088 ;
    END
  END io_rw_wdata[27]
  PIN io_rw_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.72 30.921 18.744 31.005 ;
    END
  END io_rw_wdata[28]
  PIN io_rw_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.664 0.084 17.688 ;
    END
  END io_rw_wdata[29]
  PIN io_rw_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.256 0 20.28 0.084 ;
    END
  END io_rw_wdata[2]
  PIN io_rw_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.24 0.084 18.264 ;
    END
  END io_rw_wdata[30]
  PIN io_rw_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 12.384 31.005 12.408 ;
    END
  END io_rw_wdata[31]
  PIN io_rw_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.8 0 16.824 0.084 ;
    END
  END io_rw_wdata[3]
  PIN io_rw_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.872 0 19.896 0.084 ;
    END
  END io_rw_wdata[4]
  PIN io_rw_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.728 0 13.752 0.084 ;
    END
  END io_rw_wdata[5]
  PIN io_rw_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 9.024 31.005 9.048 ;
    END
  END io_rw_wdata[6]
  PIN io_rw_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.088 0 17.112 0.084 ;
    END
  END io_rw_wdata[7]
  PIN io_rw_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.072 0 15.096 0.084 ;
    END
  END io_rw_wdata[8]
  PIN io_rw_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.784 0 14.808 0.084 ;
    END
  END io_rw_wdata[9]
  PIN io_time[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.568 0 17.592 0.084 ;
    END
  END io_time[0]
  PIN io_time[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 13.824 31.005 13.848 ;
    END
  END io_time[10]
  PIN io_time[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 12.96 31.005 12.984 ;
    END
  END io_time[11]
  PIN io_time[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 15.168 31.005 15.192 ;
    END
  END io_time[12]
  PIN io_time[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 14.496 31.005 14.52 ;
    END
  END io_time[13]
  PIN io_time[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.28 30.921 17.304 31.005 ;
    END
  END io_time[14]
  PIN io_time[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.184 30.921 17.208 31.005 ;
    END
  END io_time[15]
  PIN io_time[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.088 30.921 17.112 31.005 ;
    END
  END io_time[16]
  PIN io_time[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.144 30.921 18.168 31.005 ;
    END
  END io_time[17]
  PIN io_time[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.664 30.921 17.688 31.005 ;
    END
  END io_time[18]
  PIN io_time[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.512 30.921 16.536 31.005 ;
    END
  END io_time[19]
  PIN io_time[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.544 0 20.568 0.084 ;
    END
  END io_time[1]
  PIN io_time[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.24 30.921 18.264 31.005 ;
    END
  END io_time[20]
  PIN io_time[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.416 30.921 16.44 31.005 ;
    END
  END io_time[21]
  PIN io_time[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.224 30.921 16.248 31.005 ;
    END
  END io_time[22]
  PIN io_time[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.992 30.921 17.016 31.005 ;
    END
  END io_time[23]
  PIN io_time[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.704 30.921 16.728 31.005 ;
    END
  END io_time[24]
  PIN io_time[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.648 30.921 15.672 31.005 ;
    END
  END io_time[25]
  PIN io_time[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.032 30.921 16.056 31.005 ;
    END
  END io_time[26]
  PIN io_time[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.32 30.921 16.344 31.005 ;
    END
  END io_time[27]
  PIN io_time[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.048 30.921 18.072 31.005 ;
    END
  END io_time[28]
  PIN io_time[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.952 30.921 17.976 31.005 ;
    END
  END io_time[29]
  PIN io_time[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.352 0 20.376 0.084 ;
    END
  END io_time[2]
  PIN io_time[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.936 30.921 15.96 31.005 ;
    END
  END io_time[30]
  PIN io_time[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 11.712 31.005 11.736 ;
    END
  END io_time[31]
  PIN io_time[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.064 0 20.088 0.084 ;
    END
  END io_time[3]
  PIN io_time[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.64 0 20.664 0.084 ;
    END
  END io_time[4]
  PIN io_time[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.736 0 20.76 0.084 ;
    END
  END io_time[5]
  PIN io_time[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 9.12 31.005 9.144 ;
    END
  END io_time[6]
  PIN io_time[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 8.832 31.005 8.856 ;
    END
  END io_time[7]
  PIN io_time[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 9.984 31.005 10.008 ;
    END
  END io_time[8]
  PIN io_time[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  30.921 12.48 31.005 12.504 ;
    END
  END io_time[9]
  PIN io_tval[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.944 0.084 10.968 ;
    END
  END io_tval[0]
  PIN io_tval[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.168 0.084 15.192 ;
    END
  END io_tval[10]
  PIN io_tval[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.216 0 9.24 0.084 ;
    END
  END io_tval[11]
  PIN io_tval[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.848 0.084 10.872 ;
    END
  END io_tval[12]
  PIN io_tval[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.224 0.084 16.248 ;
    END
  END io_tval[13]
  PIN io_tval[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.76 0.084 17.784 ;
    END
  END io_tval[14]
  PIN io_tval[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.48 0 12.504 0.084 ;
    END
  END io_tval[15]
  PIN io_tval[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.144 0.084 18.168 ;
    END
  END io_tval[16]
  PIN io_tval[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.12 30.921 9.144 31.005 ;
    END
  END io_tval[17]
  PIN io_tval[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.424 0.084 23.448 ;
    END
  END io_tval[18]
  PIN io_tval[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.752 30.921 10.776 31.005 ;
    END
  END io_tval[19]
  PIN io_tval[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.928 0 8.952 0.084 ;
    END
  END io_tval[1]
  PIN io_tval[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.56 0.084 22.584 ;
    END
  END io_tval[20]
  PIN io_tval[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.04 30.921 11.064 31.005 ;
    END
  END io_tval[21]
  PIN io_tval[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.368 0.084 22.392 ;
    END
  END io_tval[22]
  PIN io_tval[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.392 30.921 7.416 31.005 ;
    END
  END io_tval[23]
  PIN io_tval[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.496 0.084 14.52 ;
    END
  END io_tval[24]
  PIN io_tval[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.504 0.084 21.528 ;
    END
  END io_tval[25]
  PIN io_tval[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  5.28 30.921 5.304 31.005 ;
    END
  END io_tval[26]
  PIN io_tval[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.352 0.084 20.376 ;
    END
  END io_tval[27]
  PIN io_tval[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.968 0.084 19.992 ;
    END
  END io_tval[28]
  PIN io_tval[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.28 0.084 17.304 ;
    END
  END io_tval[29]
  PIN io_tval[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.064 0.084 8.088 ;
    END
  END io_tval[2]
  PIN io_tval[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.912 0.084 18.936 ;
    END
  END io_tval[30]
  PIN io_tval[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.736 0 8.76 0.084 ;
    END
  END io_tval[31]
  PIN io_tval[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.64 0.084 8.664 ;
    END
  END io_tval[3]
  PIN io_tval[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.352 0.084 8.376 ;
    END
  END io_tval[4]
  PIN io_tval[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.04 0.084 11.064 ;
    END
  END io_tval[5]
  PIN io_tval[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.272 0.084 10.296 ;
    END
  END io_tval[6]
  PIN io_tval[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.52 0 11.544 0.084 ;
    END
  END io_tval[7]
  PIN io_tval[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.56 0 10.584 0.084 ;
    END
  END io_tval[8]
  PIN io_tval[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.632 0.084 13.656 ;
    END
  END io_tval[9]
  PIN io_ungated_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.504 30.921 21.528 31.005 ;
    END
  END io_ungated_clock
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.504 0 9.528 0.084 ;
    END
  END reset
  OBS
    LAYER M1 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M2 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M3 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M4 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M5 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M6 ;
     RECT  0 0 31.005 31.005 ;
    LAYER M7 ;
     RECT  0 0 31.005 31.005 ;
  END
END CSRFile
END LIBRARY
