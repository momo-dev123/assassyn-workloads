VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA run_benchmark_via1_2_57078_18_1_1585_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 1585 ;
END run_benchmark_via1_2_57078_18_1_1585_36_36

VIA run_benchmark_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END run_benchmark_VIA23_1_3_36_36

VIA run_benchmark_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END run_benchmark_VIA34_1_2_58_52

VIA run_benchmark_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END run_benchmark_VIA45_1_2_58_58

VIA run_benchmark_via5_6_120_288_1_2_58_322
  VIARULE M6_M5widePWR1p152 ;
  CUTSIZE 0.024 0.288 ;
  LAYERS M5 V5 M6 ;
  CUTSPACING 0.034 0.034 ;
  ENCLOSURE 0.019 0 0 0 ;
  ROWCOL 1 2 ;
END run_benchmark_via5_6_120_288_1_2_58_322

MACRO run_benchmark
  FOREIGN run_benchmark 0 0 ;
  CLASS BLOCK ;
  SIZE 59.121 BY 59.121 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.458 55.833 54.714 56.121 ;
        RECT  1.458 49.833 54.714 50.121 ;
        RECT  1.458 43.833 54.714 44.121 ;
        RECT  1.458 37.833 54.714 38.121 ;
        RECT  1.458 31.833 54.714 32.121 ;
        RECT  1.458 25.833 54.714 26.121 ;
        RECT  1.458 19.833 54.714 20.121 ;
        RECT  1.458 13.833 54.714 14.121 ;
        RECT  1.458 7.833 54.714 8.121 ;
        RECT  1.458 1.833 54.714 2.121 ;
      LAYER M5 ;
        RECT  54.594 1.327 54.714 58.073 ;
        RECT  48.69 1.327 48.81 58.073 ;
        RECT  42.786 1.327 42.906 58.073 ;
        RECT  36.882 1.327 37.002 58.073 ;
        RECT  30.978 1.327 31.098 58.073 ;
        RECT  25.074 1.327 25.194 58.073 ;
        RECT  19.17 1.327 19.29 58.073 ;
        RECT  13.266 1.327 13.386 58.073 ;
        RECT  7.362 1.327 7.482 58.073 ;
        RECT  1.458 1.327 1.578 58.073 ;
      LAYER M2 ;
        RECT  1.026 58.041 58.104 58.059 ;
        RECT  1.026 57.501 58.104 57.519 ;
        RECT  1.026 56.961 58.104 56.979 ;
        RECT  1.026 56.421 58.104 56.439 ;
        RECT  1.026 55.881 58.104 55.899 ;
        RECT  1.026 55.341 58.104 55.359 ;
        RECT  1.026 54.801 58.104 54.819 ;
        RECT  1.026 54.261 58.104 54.279 ;
        RECT  1.026 53.721 58.104 53.739 ;
        RECT  1.026 53.181 58.104 53.199 ;
        RECT  1.026 52.641 58.104 52.659 ;
        RECT  1.026 52.101 58.104 52.119 ;
        RECT  1.026 51.561 58.104 51.579 ;
        RECT  1.026 51.021 58.104 51.039 ;
        RECT  1.026 50.481 58.104 50.499 ;
        RECT  1.026 49.941 58.104 49.959 ;
        RECT  1.026 49.401 58.104 49.419 ;
        RECT  1.026 48.861 58.104 48.879 ;
        RECT  1.026 48.321 58.104 48.339 ;
        RECT  1.026 47.781 58.104 47.799 ;
        RECT  1.026 47.241 58.104 47.259 ;
        RECT  1.026 46.701 58.104 46.719 ;
        RECT  1.026 46.161 58.104 46.179 ;
        RECT  1.026 45.621 58.104 45.639 ;
        RECT  1.026 45.081 58.104 45.099 ;
        RECT  1.026 44.541 58.104 44.559 ;
        RECT  1.026 44.001 58.104 44.019 ;
        RECT  1.026 43.461 58.104 43.479 ;
        RECT  1.026 42.921 58.104 42.939 ;
        RECT  1.026 42.381 58.104 42.399 ;
        RECT  1.026 41.841 58.104 41.859 ;
        RECT  1.026 41.301 58.104 41.319 ;
        RECT  1.026 40.761 58.104 40.779 ;
        RECT  1.026 40.221 58.104 40.239 ;
        RECT  1.026 39.681 58.104 39.699 ;
        RECT  1.026 39.141 58.104 39.159 ;
        RECT  1.026 38.601 58.104 38.619 ;
        RECT  1.026 38.061 58.104 38.079 ;
        RECT  1.026 37.521 58.104 37.539 ;
        RECT  1.026 36.981 58.104 36.999 ;
        RECT  1.026 36.441 58.104 36.459 ;
        RECT  1.026 35.901 58.104 35.919 ;
        RECT  1.026 35.361 58.104 35.379 ;
        RECT  1.026 34.821 58.104 34.839 ;
        RECT  1.026 34.281 58.104 34.299 ;
        RECT  1.026 33.741 58.104 33.759 ;
        RECT  1.026 33.201 58.104 33.219 ;
        RECT  1.026 32.661 58.104 32.679 ;
        RECT  1.026 32.121 58.104 32.139 ;
        RECT  1.026 31.581 58.104 31.599 ;
        RECT  1.026 31.041 58.104 31.059 ;
        RECT  1.026 30.501 58.104 30.519 ;
        RECT  1.026 29.961 58.104 29.979 ;
        RECT  1.026 29.421 58.104 29.439 ;
        RECT  1.026 28.881 58.104 28.899 ;
        RECT  1.026 28.341 58.104 28.359 ;
        RECT  1.026 27.801 58.104 27.819 ;
        RECT  1.026 27.261 58.104 27.279 ;
        RECT  1.026 26.721 58.104 26.739 ;
        RECT  1.026 26.181 58.104 26.199 ;
        RECT  1.026 25.641 58.104 25.659 ;
        RECT  1.026 25.101 58.104 25.119 ;
        RECT  1.026 24.561 58.104 24.579 ;
        RECT  1.026 24.021 58.104 24.039 ;
        RECT  1.026 23.481 58.104 23.499 ;
        RECT  1.026 22.941 58.104 22.959 ;
        RECT  1.026 22.401 58.104 22.419 ;
        RECT  1.026 21.861 58.104 21.879 ;
        RECT  1.026 21.321 58.104 21.339 ;
        RECT  1.026 20.781 58.104 20.799 ;
        RECT  1.026 20.241 58.104 20.259 ;
        RECT  1.026 19.701 58.104 19.719 ;
        RECT  1.026 19.161 58.104 19.179 ;
        RECT  1.026 18.621 58.104 18.639 ;
        RECT  1.026 18.081 58.104 18.099 ;
        RECT  1.026 17.541 58.104 17.559 ;
        RECT  1.026 17.001 58.104 17.019 ;
        RECT  1.026 16.461 58.104 16.479 ;
        RECT  1.026 15.921 58.104 15.939 ;
        RECT  1.026 15.381 58.104 15.399 ;
        RECT  1.026 14.841 58.104 14.859 ;
        RECT  1.026 14.301 58.104 14.319 ;
        RECT  1.026 13.761 58.104 13.779 ;
        RECT  1.026 13.221 58.104 13.239 ;
        RECT  1.026 12.681 58.104 12.699 ;
        RECT  1.026 12.141 58.104 12.159 ;
        RECT  1.026 11.601 58.104 11.619 ;
        RECT  1.026 11.061 58.104 11.079 ;
        RECT  1.026 10.521 58.104 10.539 ;
        RECT  1.026 9.981 58.104 9.999 ;
        RECT  1.026 9.441 58.104 9.459 ;
        RECT  1.026 8.901 58.104 8.919 ;
        RECT  1.026 8.361 58.104 8.379 ;
        RECT  1.026 7.821 58.104 7.839 ;
        RECT  1.026 7.281 58.104 7.299 ;
        RECT  1.026 6.741 58.104 6.759 ;
        RECT  1.026 6.201 58.104 6.219 ;
        RECT  1.026 5.661 58.104 5.679 ;
        RECT  1.026 5.121 58.104 5.139 ;
        RECT  1.026 4.581 58.104 4.599 ;
        RECT  1.026 4.041 58.104 4.059 ;
        RECT  1.026 3.501 58.104 3.519 ;
        RECT  1.026 2.961 58.104 2.979 ;
        RECT  1.026 2.421 58.104 2.439 ;
        RECT  1.026 1.881 58.104 1.899 ;
        RECT  1.026 1.341 58.104 1.359 ;
      LAYER M1 ;
        RECT  1.026 58.041 58.104 58.059 ;
        RECT  1.026 57.501 58.104 57.519 ;
        RECT  1.026 56.961 58.104 56.979 ;
        RECT  1.026 56.421 58.104 56.439 ;
        RECT  1.026 55.881 58.104 55.899 ;
        RECT  1.026 55.341 58.104 55.359 ;
        RECT  1.026 54.801 58.104 54.819 ;
        RECT  1.026 54.261 58.104 54.279 ;
        RECT  1.026 53.721 58.104 53.739 ;
        RECT  1.026 53.181 58.104 53.199 ;
        RECT  1.026 52.641 58.104 52.659 ;
        RECT  1.026 52.101 58.104 52.119 ;
        RECT  1.026 51.561 58.104 51.579 ;
        RECT  1.026 51.021 58.104 51.039 ;
        RECT  1.026 50.481 58.104 50.499 ;
        RECT  1.026 49.941 58.104 49.959 ;
        RECT  1.026 49.401 58.104 49.419 ;
        RECT  1.026 48.861 58.104 48.879 ;
        RECT  1.026 48.321 58.104 48.339 ;
        RECT  1.026 47.781 58.104 47.799 ;
        RECT  1.026 47.241 58.104 47.259 ;
        RECT  1.026 46.701 58.104 46.719 ;
        RECT  1.026 46.161 58.104 46.179 ;
        RECT  1.026 45.621 58.104 45.639 ;
        RECT  1.026 45.081 58.104 45.099 ;
        RECT  1.026 44.541 58.104 44.559 ;
        RECT  1.026 44.001 58.104 44.019 ;
        RECT  1.026 43.461 58.104 43.479 ;
        RECT  1.026 42.921 58.104 42.939 ;
        RECT  1.026 42.381 58.104 42.399 ;
        RECT  1.026 41.841 58.104 41.859 ;
        RECT  1.026 41.301 58.104 41.319 ;
        RECT  1.026 40.761 58.104 40.779 ;
        RECT  1.026 40.221 58.104 40.239 ;
        RECT  1.026 39.681 58.104 39.699 ;
        RECT  1.026 39.141 58.104 39.159 ;
        RECT  1.026 38.601 58.104 38.619 ;
        RECT  1.026 38.061 58.104 38.079 ;
        RECT  1.026 37.521 58.104 37.539 ;
        RECT  1.026 36.981 58.104 36.999 ;
        RECT  1.026 36.441 58.104 36.459 ;
        RECT  1.026 35.901 58.104 35.919 ;
        RECT  1.026 35.361 58.104 35.379 ;
        RECT  1.026 34.821 58.104 34.839 ;
        RECT  1.026 34.281 58.104 34.299 ;
        RECT  1.026 33.741 58.104 33.759 ;
        RECT  1.026 33.201 58.104 33.219 ;
        RECT  1.026 32.661 58.104 32.679 ;
        RECT  1.026 32.121 58.104 32.139 ;
        RECT  1.026 31.581 58.104 31.599 ;
        RECT  1.026 31.041 58.104 31.059 ;
        RECT  1.026 30.501 58.104 30.519 ;
        RECT  1.026 29.961 58.104 29.979 ;
        RECT  1.026 29.421 58.104 29.439 ;
        RECT  1.026 28.881 58.104 28.899 ;
        RECT  1.026 28.341 58.104 28.359 ;
        RECT  1.026 27.801 58.104 27.819 ;
        RECT  1.026 27.261 58.104 27.279 ;
        RECT  1.026 26.721 58.104 26.739 ;
        RECT  1.026 26.181 58.104 26.199 ;
        RECT  1.026 25.641 58.104 25.659 ;
        RECT  1.026 25.101 58.104 25.119 ;
        RECT  1.026 24.561 58.104 24.579 ;
        RECT  1.026 24.021 58.104 24.039 ;
        RECT  1.026 23.481 58.104 23.499 ;
        RECT  1.026 22.941 58.104 22.959 ;
        RECT  1.026 22.401 58.104 22.419 ;
        RECT  1.026 21.861 58.104 21.879 ;
        RECT  1.026 21.321 58.104 21.339 ;
        RECT  1.026 20.781 58.104 20.799 ;
        RECT  1.026 20.241 58.104 20.259 ;
        RECT  1.026 19.701 58.104 19.719 ;
        RECT  1.026 19.161 58.104 19.179 ;
        RECT  1.026 18.621 58.104 18.639 ;
        RECT  1.026 18.081 58.104 18.099 ;
        RECT  1.026 17.541 58.104 17.559 ;
        RECT  1.026 17.001 58.104 17.019 ;
        RECT  1.026 16.461 58.104 16.479 ;
        RECT  1.026 15.921 58.104 15.939 ;
        RECT  1.026 15.381 58.104 15.399 ;
        RECT  1.026 14.841 58.104 14.859 ;
        RECT  1.026 14.301 58.104 14.319 ;
        RECT  1.026 13.761 58.104 13.779 ;
        RECT  1.026 13.221 58.104 13.239 ;
        RECT  1.026 12.681 58.104 12.699 ;
        RECT  1.026 12.141 58.104 12.159 ;
        RECT  1.026 11.601 58.104 11.619 ;
        RECT  1.026 11.061 58.104 11.079 ;
        RECT  1.026 10.521 58.104 10.539 ;
        RECT  1.026 9.981 58.104 9.999 ;
        RECT  1.026 9.441 58.104 9.459 ;
        RECT  1.026 8.901 58.104 8.919 ;
        RECT  1.026 8.361 58.104 8.379 ;
        RECT  1.026 7.821 58.104 7.839 ;
        RECT  1.026 7.281 58.104 7.299 ;
        RECT  1.026 6.741 58.104 6.759 ;
        RECT  1.026 6.201 58.104 6.219 ;
        RECT  1.026 5.661 58.104 5.679 ;
        RECT  1.026 5.121 58.104 5.139 ;
        RECT  1.026 4.581 58.104 4.599 ;
        RECT  1.026 4.041 58.104 4.059 ;
        RECT  1.026 3.501 58.104 3.519 ;
        RECT  1.026 2.961 58.104 2.979 ;
        RECT  1.026 2.421 58.104 2.439 ;
        RECT  1.026 1.881 58.104 1.899 ;
        RECT  1.026 1.341 58.104 1.359 ;
      VIA 54.654 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.75 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.846 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 55.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 49.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 43.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.654 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 58.033 54.699 58.067 ;
      VIA 54.654 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 57.493 54.699 57.527 ;
      VIA 54.654 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 56.953 54.699 56.987 ;
      VIA 54.654 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 56.413 54.699 56.447 ;
      VIA 54.654 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 55.873 54.699 55.907 ;
      VIA 54.654 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 55.333 54.699 55.367 ;
      VIA 54.654 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 54.793 54.699 54.827 ;
      VIA 54.654 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 54.253 54.699 54.287 ;
      VIA 54.654 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 53.713 54.699 53.747 ;
      VIA 54.654 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 53.173 54.699 53.207 ;
      VIA 54.654 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 52.633 54.699 52.667 ;
      VIA 54.654 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 52.093 54.699 52.127 ;
      VIA 54.654 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 51.553 54.699 51.587 ;
      VIA 54.654 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 51.013 54.699 51.047 ;
      VIA 54.654 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 50.473 54.699 50.507 ;
      VIA 54.654 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 49.933 54.699 49.967 ;
      VIA 54.654 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 49.393 54.699 49.427 ;
      VIA 54.654 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 48.853 54.699 48.887 ;
      VIA 54.654 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 48.313 54.699 48.347 ;
      VIA 54.654 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 47.773 54.699 47.807 ;
      VIA 54.654 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 47.233 54.699 47.267 ;
      VIA 54.654 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 46.693 54.699 46.727 ;
      VIA 54.654 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 46.153 54.699 46.187 ;
      VIA 54.654 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 45.613 54.699 45.647 ;
      VIA 54.654 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 45.073 54.699 45.107 ;
      VIA 54.654 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 44.533 54.699 44.567 ;
      VIA 54.654 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 43.993 54.699 44.027 ;
      VIA 54.654 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 43.453 54.699 43.487 ;
      VIA 54.654 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 42.913 54.699 42.947 ;
      VIA 54.654 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 42.373 54.699 42.407 ;
      VIA 54.654 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 41.833 54.699 41.867 ;
      VIA 54.654 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 41.293 54.699 41.327 ;
      VIA 54.654 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 40.753 54.699 40.787 ;
      VIA 54.654 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 40.213 54.699 40.247 ;
      VIA 54.654 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 39.673 54.699 39.707 ;
      VIA 54.654 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 39.133 54.699 39.167 ;
      VIA 54.654 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 38.593 54.699 38.627 ;
      VIA 54.654 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 38.053 54.699 38.087 ;
      VIA 54.654 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 37.513 54.699 37.547 ;
      VIA 54.654 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 36.973 54.699 37.007 ;
      VIA 54.654 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 36.433 54.699 36.467 ;
      VIA 54.654 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 35.893 54.699 35.927 ;
      VIA 54.654 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 35.353 54.699 35.387 ;
      VIA 54.654 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 34.813 54.699 34.847 ;
      VIA 54.654 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 34.273 54.699 34.307 ;
      VIA 54.654 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 33.733 54.699 33.767 ;
      VIA 54.654 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 33.193 54.699 33.227 ;
      VIA 54.654 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 32.653 54.699 32.687 ;
      VIA 54.654 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 32.113 54.699 32.147 ;
      VIA 54.654 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 31.573 54.699 31.607 ;
      VIA 54.654 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 31.033 54.699 31.067 ;
      VIA 54.654 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 30.493 54.699 30.527 ;
      VIA 54.654 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 29.953 54.699 29.987 ;
      VIA 54.654 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 29.413 54.699 29.447 ;
      VIA 54.654 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 28.873 54.699 28.907 ;
      VIA 54.654 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 28.333 54.699 28.367 ;
      VIA 54.654 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 27.793 54.699 27.827 ;
      VIA 54.654 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 27.253 54.699 27.287 ;
      VIA 54.654 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 26.713 54.699 26.747 ;
      VIA 54.654 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 26.173 54.699 26.207 ;
      VIA 54.654 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 25.633 54.699 25.667 ;
      VIA 54.654 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 25.093 54.699 25.127 ;
      VIA 54.654 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 24.553 54.699 24.587 ;
      VIA 54.654 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 24.013 54.699 24.047 ;
      VIA 54.654 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 23.473 54.699 23.507 ;
      VIA 54.654 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 22.933 54.699 22.967 ;
      VIA 54.654 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 22.393 54.699 22.427 ;
      VIA 54.654 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 21.853 54.699 21.887 ;
      VIA 54.654 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 21.313 54.699 21.347 ;
      VIA 54.654 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 20.773 54.699 20.807 ;
      VIA 54.654 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 20.233 54.699 20.267 ;
      VIA 54.654 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 19.693 54.699 19.727 ;
      VIA 54.654 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 19.153 54.699 19.187 ;
      VIA 54.654 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 18.613 54.699 18.647 ;
      VIA 54.654 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 18.073 54.699 18.107 ;
      VIA 54.654 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 17.533 54.699 17.567 ;
      VIA 54.654 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 16.993 54.699 17.027 ;
      VIA 54.654 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 16.453 54.699 16.487 ;
      VIA 54.654 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 15.913 54.699 15.947 ;
      VIA 54.654 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 15.373 54.699 15.407 ;
      VIA 54.654 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 14.833 54.699 14.867 ;
      VIA 54.654 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 14.293 54.699 14.327 ;
      VIA 54.654 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 13.753 54.699 13.787 ;
      VIA 54.654 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 13.213 54.699 13.247 ;
      VIA 54.654 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 12.673 54.699 12.707 ;
      VIA 54.654 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 12.133 54.699 12.167 ;
      VIA 54.654 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 11.593 54.699 11.627 ;
      VIA 54.654 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 11.053 54.699 11.087 ;
      VIA 54.654 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 10.513 54.699 10.547 ;
      VIA 54.654 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 9.973 54.699 10.007 ;
      VIA 54.654 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 9.433 54.699 9.467 ;
      VIA 54.654 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 8.893 54.699 8.927 ;
      VIA 54.654 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 8.353 54.699 8.387 ;
      VIA 54.654 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 7.813 54.699 7.847 ;
      VIA 54.654 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 7.273 54.699 7.307 ;
      VIA 54.654 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 6.733 54.699 6.767 ;
      VIA 54.654 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 6.193 54.699 6.227 ;
      VIA 54.654 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 5.653 54.699 5.687 ;
      VIA 54.654 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 5.113 54.699 5.147 ;
      VIA 54.654 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 4.573 54.699 4.607 ;
      VIA 54.654 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 4.033 54.699 4.067 ;
      VIA 54.654 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 3.493 54.699 3.527 ;
      VIA 54.654 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 2.953 54.699 2.987 ;
      VIA 54.654 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 2.413 54.699 2.447 ;
      VIA 54.654 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 1.873 54.699 1.907 ;
      VIA 54.654 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.654 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.609 1.333 54.699 1.367 ;
      VIA 54.654 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.654 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 58.033 48.795 58.067 ;
      VIA 48.75 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 57.493 48.795 57.527 ;
      VIA 48.75 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 56.953 48.795 56.987 ;
      VIA 48.75 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 56.413 48.795 56.447 ;
      VIA 48.75 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 55.873 48.795 55.907 ;
      VIA 48.75 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 55.333 48.795 55.367 ;
      VIA 48.75 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 54.793 48.795 54.827 ;
      VIA 48.75 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 54.253 48.795 54.287 ;
      VIA 48.75 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 53.713 48.795 53.747 ;
      VIA 48.75 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 53.173 48.795 53.207 ;
      VIA 48.75 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 52.633 48.795 52.667 ;
      VIA 48.75 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 52.093 48.795 52.127 ;
      VIA 48.75 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 51.553 48.795 51.587 ;
      VIA 48.75 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 51.013 48.795 51.047 ;
      VIA 48.75 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 50.473 48.795 50.507 ;
      VIA 48.75 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 49.933 48.795 49.967 ;
      VIA 48.75 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 49.393 48.795 49.427 ;
      VIA 48.75 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 48.853 48.795 48.887 ;
      VIA 48.75 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 48.313 48.795 48.347 ;
      VIA 48.75 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 47.773 48.795 47.807 ;
      VIA 48.75 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 47.233 48.795 47.267 ;
      VIA 48.75 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 46.693 48.795 46.727 ;
      VIA 48.75 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 46.153 48.795 46.187 ;
      VIA 48.75 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 45.613 48.795 45.647 ;
      VIA 48.75 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 45.073 48.795 45.107 ;
      VIA 48.75 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 44.533 48.795 44.567 ;
      VIA 48.75 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 43.993 48.795 44.027 ;
      VIA 48.75 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 43.453 48.795 43.487 ;
      VIA 48.75 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 42.913 48.795 42.947 ;
      VIA 48.75 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 42.373 48.795 42.407 ;
      VIA 48.75 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 41.833 48.795 41.867 ;
      VIA 48.75 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 41.293 48.795 41.327 ;
      VIA 48.75 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 40.753 48.795 40.787 ;
      VIA 48.75 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 40.213 48.795 40.247 ;
      VIA 48.75 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 39.673 48.795 39.707 ;
      VIA 48.75 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 39.133 48.795 39.167 ;
      VIA 48.75 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 38.593 48.795 38.627 ;
      VIA 48.75 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 38.053 48.795 38.087 ;
      VIA 48.75 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 37.513 48.795 37.547 ;
      VIA 48.75 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 36.973 48.795 37.007 ;
      VIA 48.75 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 36.433 48.795 36.467 ;
      VIA 48.75 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 35.893 48.795 35.927 ;
      VIA 48.75 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 35.353 48.795 35.387 ;
      VIA 48.75 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 34.813 48.795 34.847 ;
      VIA 48.75 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 34.273 48.795 34.307 ;
      VIA 48.75 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 33.733 48.795 33.767 ;
      VIA 48.75 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 33.193 48.795 33.227 ;
      VIA 48.75 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 32.653 48.795 32.687 ;
      VIA 48.75 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 32.113 48.795 32.147 ;
      VIA 48.75 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 31.573 48.795 31.607 ;
      VIA 48.75 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 31.033 48.795 31.067 ;
      VIA 48.75 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 30.493 48.795 30.527 ;
      VIA 48.75 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 29.953 48.795 29.987 ;
      VIA 48.75 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 29.413 48.795 29.447 ;
      VIA 48.75 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 28.873 48.795 28.907 ;
      VIA 48.75 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 28.333 48.795 28.367 ;
      VIA 48.75 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 27.793 48.795 27.827 ;
      VIA 48.75 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 27.253 48.795 27.287 ;
      VIA 48.75 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 26.713 48.795 26.747 ;
      VIA 48.75 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 26.173 48.795 26.207 ;
      VIA 48.75 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 25.633 48.795 25.667 ;
      VIA 48.75 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 25.093 48.795 25.127 ;
      VIA 48.75 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 24.553 48.795 24.587 ;
      VIA 48.75 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 24.013 48.795 24.047 ;
      VIA 48.75 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 23.473 48.795 23.507 ;
      VIA 48.75 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 22.933 48.795 22.967 ;
      VIA 48.75 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 22.393 48.795 22.427 ;
      VIA 48.75 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 21.853 48.795 21.887 ;
      VIA 48.75 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 21.313 48.795 21.347 ;
      VIA 48.75 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 20.773 48.795 20.807 ;
      VIA 48.75 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 20.233 48.795 20.267 ;
      VIA 48.75 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 19.693 48.795 19.727 ;
      VIA 48.75 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 19.153 48.795 19.187 ;
      VIA 48.75 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 18.613 48.795 18.647 ;
      VIA 48.75 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 18.073 48.795 18.107 ;
      VIA 48.75 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 17.533 48.795 17.567 ;
      VIA 48.75 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 16.993 48.795 17.027 ;
      VIA 48.75 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 16.453 48.795 16.487 ;
      VIA 48.75 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 15.913 48.795 15.947 ;
      VIA 48.75 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 15.373 48.795 15.407 ;
      VIA 48.75 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 14.833 48.795 14.867 ;
      VIA 48.75 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 14.293 48.795 14.327 ;
      VIA 48.75 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 13.753 48.795 13.787 ;
      VIA 48.75 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 13.213 48.795 13.247 ;
      VIA 48.75 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 12.673 48.795 12.707 ;
      VIA 48.75 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 12.133 48.795 12.167 ;
      VIA 48.75 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 11.593 48.795 11.627 ;
      VIA 48.75 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 11.053 48.795 11.087 ;
      VIA 48.75 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 10.513 48.795 10.547 ;
      VIA 48.75 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 9.973 48.795 10.007 ;
      VIA 48.75 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 9.433 48.795 9.467 ;
      VIA 48.75 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 8.893 48.795 8.927 ;
      VIA 48.75 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 8.353 48.795 8.387 ;
      VIA 48.75 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 7.813 48.795 7.847 ;
      VIA 48.75 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 7.273 48.795 7.307 ;
      VIA 48.75 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 6.733 48.795 6.767 ;
      VIA 48.75 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 6.193 48.795 6.227 ;
      VIA 48.75 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 5.653 48.795 5.687 ;
      VIA 48.75 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 5.113 48.795 5.147 ;
      VIA 48.75 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 4.573 48.795 4.607 ;
      VIA 48.75 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 4.033 48.795 4.067 ;
      VIA 48.75 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 3.493 48.795 3.527 ;
      VIA 48.75 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 2.953 48.795 2.987 ;
      VIA 48.75 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 2.413 48.795 2.447 ;
      VIA 48.75 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 1.873 48.795 1.907 ;
      VIA 48.75 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.75 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.705 1.333 48.795 1.367 ;
      VIA 48.75 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.75 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 58.033 42.891 58.067 ;
      VIA 42.846 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 57.493 42.891 57.527 ;
      VIA 42.846 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 56.953 42.891 56.987 ;
      VIA 42.846 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 56.413 42.891 56.447 ;
      VIA 42.846 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 55.873 42.891 55.907 ;
      VIA 42.846 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 55.333 42.891 55.367 ;
      VIA 42.846 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 54.793 42.891 54.827 ;
      VIA 42.846 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 54.253 42.891 54.287 ;
      VIA 42.846 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 53.713 42.891 53.747 ;
      VIA 42.846 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 53.173 42.891 53.207 ;
      VIA 42.846 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 52.633 42.891 52.667 ;
      VIA 42.846 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 52.093 42.891 52.127 ;
      VIA 42.846 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 51.553 42.891 51.587 ;
      VIA 42.846 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 51.013 42.891 51.047 ;
      VIA 42.846 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 50.473 42.891 50.507 ;
      VIA 42.846 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 49.933 42.891 49.967 ;
      VIA 42.846 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 49.393 42.891 49.427 ;
      VIA 42.846 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 48.853 42.891 48.887 ;
      VIA 42.846 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 48.313 42.891 48.347 ;
      VIA 42.846 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 47.773 42.891 47.807 ;
      VIA 42.846 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 47.233 42.891 47.267 ;
      VIA 42.846 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 46.693 42.891 46.727 ;
      VIA 42.846 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 46.153 42.891 46.187 ;
      VIA 42.846 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 45.613 42.891 45.647 ;
      VIA 42.846 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 45.073 42.891 45.107 ;
      VIA 42.846 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 44.533 42.891 44.567 ;
      VIA 42.846 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 43.993 42.891 44.027 ;
      VIA 42.846 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 43.453 42.891 43.487 ;
      VIA 42.846 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 42.913 42.891 42.947 ;
      VIA 42.846 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 42.373 42.891 42.407 ;
      VIA 42.846 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 41.833 42.891 41.867 ;
      VIA 42.846 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 41.293 42.891 41.327 ;
      VIA 42.846 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 40.753 42.891 40.787 ;
      VIA 42.846 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 40.213 42.891 40.247 ;
      VIA 42.846 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 39.673 42.891 39.707 ;
      VIA 42.846 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 39.133 42.891 39.167 ;
      VIA 42.846 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 38.593 42.891 38.627 ;
      VIA 42.846 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 38.053 42.891 38.087 ;
      VIA 42.846 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 37.513 42.891 37.547 ;
      VIA 42.846 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 36.973 42.891 37.007 ;
      VIA 42.846 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 36.433 42.891 36.467 ;
      VIA 42.846 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 35.893 42.891 35.927 ;
      VIA 42.846 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 35.353 42.891 35.387 ;
      VIA 42.846 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 34.813 42.891 34.847 ;
      VIA 42.846 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 34.273 42.891 34.307 ;
      VIA 42.846 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 33.733 42.891 33.767 ;
      VIA 42.846 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 33.193 42.891 33.227 ;
      VIA 42.846 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 32.653 42.891 32.687 ;
      VIA 42.846 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 32.113 42.891 32.147 ;
      VIA 42.846 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 31.573 42.891 31.607 ;
      VIA 42.846 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 31.033 42.891 31.067 ;
      VIA 42.846 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 30.493 42.891 30.527 ;
      VIA 42.846 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 29.953 42.891 29.987 ;
      VIA 42.846 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 29.413 42.891 29.447 ;
      VIA 42.846 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 28.873 42.891 28.907 ;
      VIA 42.846 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 28.333 42.891 28.367 ;
      VIA 42.846 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 27.793 42.891 27.827 ;
      VIA 42.846 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 27.253 42.891 27.287 ;
      VIA 42.846 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 26.713 42.891 26.747 ;
      VIA 42.846 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 26.173 42.891 26.207 ;
      VIA 42.846 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 25.633 42.891 25.667 ;
      VIA 42.846 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 25.093 42.891 25.127 ;
      VIA 42.846 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 24.553 42.891 24.587 ;
      VIA 42.846 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 24.013 42.891 24.047 ;
      VIA 42.846 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 23.473 42.891 23.507 ;
      VIA 42.846 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 22.933 42.891 22.967 ;
      VIA 42.846 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 22.393 42.891 22.427 ;
      VIA 42.846 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 21.853 42.891 21.887 ;
      VIA 42.846 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 21.313 42.891 21.347 ;
      VIA 42.846 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 20.773 42.891 20.807 ;
      VIA 42.846 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 20.233 42.891 20.267 ;
      VIA 42.846 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 19.693 42.891 19.727 ;
      VIA 42.846 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 19.153 42.891 19.187 ;
      VIA 42.846 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 18.613 42.891 18.647 ;
      VIA 42.846 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 18.073 42.891 18.107 ;
      VIA 42.846 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 17.533 42.891 17.567 ;
      VIA 42.846 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 16.993 42.891 17.027 ;
      VIA 42.846 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 16.453 42.891 16.487 ;
      VIA 42.846 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 15.913 42.891 15.947 ;
      VIA 42.846 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 15.373 42.891 15.407 ;
      VIA 42.846 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 14.833 42.891 14.867 ;
      VIA 42.846 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 14.293 42.891 14.327 ;
      VIA 42.846 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 13.753 42.891 13.787 ;
      VIA 42.846 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 13.213 42.891 13.247 ;
      VIA 42.846 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 12.673 42.891 12.707 ;
      VIA 42.846 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 12.133 42.891 12.167 ;
      VIA 42.846 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 11.593 42.891 11.627 ;
      VIA 42.846 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 11.053 42.891 11.087 ;
      VIA 42.846 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 10.513 42.891 10.547 ;
      VIA 42.846 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 9.973 42.891 10.007 ;
      VIA 42.846 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 9.433 42.891 9.467 ;
      VIA 42.846 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 8.893 42.891 8.927 ;
      VIA 42.846 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 8.353 42.891 8.387 ;
      VIA 42.846 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 7.813 42.891 7.847 ;
      VIA 42.846 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 7.273 42.891 7.307 ;
      VIA 42.846 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 6.733 42.891 6.767 ;
      VIA 42.846 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 6.193 42.891 6.227 ;
      VIA 42.846 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 5.653 42.891 5.687 ;
      VIA 42.846 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 5.113 42.891 5.147 ;
      VIA 42.846 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 4.573 42.891 4.607 ;
      VIA 42.846 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 4.033 42.891 4.067 ;
      VIA 42.846 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 3.493 42.891 3.527 ;
      VIA 42.846 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 2.953 42.891 2.987 ;
      VIA 42.846 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 2.413 42.891 2.447 ;
      VIA 42.846 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 1.873 42.891 1.907 ;
      VIA 42.846 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.846 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.801 1.333 42.891 1.367 ;
      VIA 42.846 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.846 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 58.033 36.987 58.067 ;
      VIA 36.942 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 57.493 36.987 57.527 ;
      VIA 36.942 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 56.953 36.987 56.987 ;
      VIA 36.942 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 56.413 36.987 56.447 ;
      VIA 36.942 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 55.873 36.987 55.907 ;
      VIA 36.942 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 55.333 36.987 55.367 ;
      VIA 36.942 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 54.793 36.987 54.827 ;
      VIA 36.942 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 54.253 36.987 54.287 ;
      VIA 36.942 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 53.713 36.987 53.747 ;
      VIA 36.942 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 53.173 36.987 53.207 ;
      VIA 36.942 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 52.633 36.987 52.667 ;
      VIA 36.942 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 52.093 36.987 52.127 ;
      VIA 36.942 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 51.553 36.987 51.587 ;
      VIA 36.942 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 51.013 36.987 51.047 ;
      VIA 36.942 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 50.473 36.987 50.507 ;
      VIA 36.942 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 49.933 36.987 49.967 ;
      VIA 36.942 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 49.393 36.987 49.427 ;
      VIA 36.942 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 48.853 36.987 48.887 ;
      VIA 36.942 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 48.313 36.987 48.347 ;
      VIA 36.942 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 47.773 36.987 47.807 ;
      VIA 36.942 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 47.233 36.987 47.267 ;
      VIA 36.942 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 46.693 36.987 46.727 ;
      VIA 36.942 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 46.153 36.987 46.187 ;
      VIA 36.942 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 45.613 36.987 45.647 ;
      VIA 36.942 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 45.073 36.987 45.107 ;
      VIA 36.942 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 44.533 36.987 44.567 ;
      VIA 36.942 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 43.993 36.987 44.027 ;
      VIA 36.942 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 43.453 36.987 43.487 ;
      VIA 36.942 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 42.913 36.987 42.947 ;
      VIA 36.942 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 42.373 36.987 42.407 ;
      VIA 36.942 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 41.833 36.987 41.867 ;
      VIA 36.942 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 41.293 36.987 41.327 ;
      VIA 36.942 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 40.753 36.987 40.787 ;
      VIA 36.942 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 40.213 36.987 40.247 ;
      VIA 36.942 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.673 36.987 39.707 ;
      VIA 36.942 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.133 36.987 39.167 ;
      VIA 36.942 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.593 36.987 38.627 ;
      VIA 36.942 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.053 36.987 38.087 ;
      VIA 36.942 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 37.513 36.987 37.547 ;
      VIA 36.942 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.973 36.987 37.007 ;
      VIA 36.942 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.433 36.987 36.467 ;
      VIA 36.942 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.893 36.987 35.927 ;
      VIA 36.942 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.353 36.987 35.387 ;
      VIA 36.942 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.813 36.987 34.847 ;
      VIA 36.942 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.273 36.987 34.307 ;
      VIA 36.942 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.733 36.987 33.767 ;
      VIA 36.942 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.193 36.987 33.227 ;
      VIA 36.942 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.653 36.987 32.687 ;
      VIA 36.942 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.113 36.987 32.147 ;
      VIA 36.942 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.573 36.987 31.607 ;
      VIA 36.942 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.033 36.987 31.067 ;
      VIA 36.942 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 30.493 36.987 30.527 ;
      VIA 36.942 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.953 36.987 29.987 ;
      VIA 36.942 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.413 36.987 29.447 ;
      VIA 36.942 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.873 36.987 28.907 ;
      VIA 36.942 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.333 36.987 28.367 ;
      VIA 36.942 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.793 36.987 27.827 ;
      VIA 36.942 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.253 36.987 27.287 ;
      VIA 36.942 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.713 36.987 26.747 ;
      VIA 36.942 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.173 36.987 26.207 ;
      VIA 36.942 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.633 36.987 25.667 ;
      VIA 36.942 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.093 36.987 25.127 ;
      VIA 36.942 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.553 36.987 24.587 ;
      VIA 36.942 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.013 36.987 24.047 ;
      VIA 36.942 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 23.473 36.987 23.507 ;
      VIA 36.942 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.933 36.987 22.967 ;
      VIA 36.942 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.393 36.987 22.427 ;
      VIA 36.942 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.853 36.987 21.887 ;
      VIA 36.942 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.313 36.987 21.347 ;
      VIA 36.942 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.773 36.987 20.807 ;
      VIA 36.942 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.233 36.987 20.267 ;
      VIA 36.942 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.693 36.987 19.727 ;
      VIA 36.942 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.153 36.987 19.187 ;
      VIA 36.942 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.613 36.987 18.647 ;
      VIA 36.942 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.073 36.987 18.107 ;
      VIA 36.942 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 17.533 36.987 17.567 ;
      VIA 36.942 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.993 36.987 17.027 ;
      VIA 36.942 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.453 36.987 16.487 ;
      VIA 36.942 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.913 36.987 15.947 ;
      VIA 36.942 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.373 36.987 15.407 ;
      VIA 36.942 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.833 36.987 14.867 ;
      VIA 36.942 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.293 36.987 14.327 ;
      VIA 36.942 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.753 36.987 13.787 ;
      VIA 36.942 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.213 36.987 13.247 ;
      VIA 36.942 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.673 36.987 12.707 ;
      VIA 36.942 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.133 36.987 12.167 ;
      VIA 36.942 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.593 36.987 11.627 ;
      VIA 36.942 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.053 36.987 11.087 ;
      VIA 36.942 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 10.513 36.987 10.547 ;
      VIA 36.942 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.973 36.987 10.007 ;
      VIA 36.942 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.433 36.987 9.467 ;
      VIA 36.942 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.893 36.987 8.927 ;
      VIA 36.942 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.353 36.987 8.387 ;
      VIA 36.942 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.813 36.987 7.847 ;
      VIA 36.942 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.273 36.987 7.307 ;
      VIA 36.942 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.733 36.987 6.767 ;
      VIA 36.942 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.193 36.987 6.227 ;
      VIA 36.942 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.653 36.987 5.687 ;
      VIA 36.942 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.113 36.987 5.147 ;
      VIA 36.942 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.573 36.987 4.607 ;
      VIA 36.942 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.033 36.987 4.067 ;
      VIA 36.942 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 3.493 36.987 3.527 ;
      VIA 36.942 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.953 36.987 2.987 ;
      VIA 36.942 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.413 36.987 2.447 ;
      VIA 36.942 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.873 36.987 1.907 ;
      VIA 36.942 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.333 36.987 1.367 ;
      VIA 36.942 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 58.033 31.083 58.067 ;
      VIA 31.038 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 57.493 31.083 57.527 ;
      VIA 31.038 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 56.953 31.083 56.987 ;
      VIA 31.038 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 56.413 31.083 56.447 ;
      VIA 31.038 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 55.873 31.083 55.907 ;
      VIA 31.038 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 55.333 31.083 55.367 ;
      VIA 31.038 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 54.793 31.083 54.827 ;
      VIA 31.038 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 54.253 31.083 54.287 ;
      VIA 31.038 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 53.713 31.083 53.747 ;
      VIA 31.038 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 53.173 31.083 53.207 ;
      VIA 31.038 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 52.633 31.083 52.667 ;
      VIA 31.038 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 52.093 31.083 52.127 ;
      VIA 31.038 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 51.553 31.083 51.587 ;
      VIA 31.038 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 51.013 31.083 51.047 ;
      VIA 31.038 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 50.473 31.083 50.507 ;
      VIA 31.038 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 49.933 31.083 49.967 ;
      VIA 31.038 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 49.393 31.083 49.427 ;
      VIA 31.038 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 48.853 31.083 48.887 ;
      VIA 31.038 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 48.313 31.083 48.347 ;
      VIA 31.038 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 47.773 31.083 47.807 ;
      VIA 31.038 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 47.233 31.083 47.267 ;
      VIA 31.038 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 46.693 31.083 46.727 ;
      VIA 31.038 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 46.153 31.083 46.187 ;
      VIA 31.038 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 45.613 31.083 45.647 ;
      VIA 31.038 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 45.073 31.083 45.107 ;
      VIA 31.038 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 44.533 31.083 44.567 ;
      VIA 31.038 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 43.993 31.083 44.027 ;
      VIA 31.038 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 43.453 31.083 43.487 ;
      VIA 31.038 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 42.913 31.083 42.947 ;
      VIA 31.038 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 42.373 31.083 42.407 ;
      VIA 31.038 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 41.833 31.083 41.867 ;
      VIA 31.038 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 41.293 31.083 41.327 ;
      VIA 31.038 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 40.753 31.083 40.787 ;
      VIA 31.038 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 40.213 31.083 40.247 ;
      VIA 31.038 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.673 31.083 39.707 ;
      VIA 31.038 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.133 31.083 39.167 ;
      VIA 31.038 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.593 31.083 38.627 ;
      VIA 31.038 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.053 31.083 38.087 ;
      VIA 31.038 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 37.513 31.083 37.547 ;
      VIA 31.038 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.973 31.083 37.007 ;
      VIA 31.038 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.433 31.083 36.467 ;
      VIA 31.038 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.893 31.083 35.927 ;
      VIA 31.038 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.353 31.083 35.387 ;
      VIA 31.038 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.813 31.083 34.847 ;
      VIA 31.038 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.273 31.083 34.307 ;
      VIA 31.038 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.733 31.083 33.767 ;
      VIA 31.038 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.193 31.083 33.227 ;
      VIA 31.038 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.653 31.083 32.687 ;
      VIA 31.038 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.113 31.083 32.147 ;
      VIA 31.038 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.573 31.083 31.607 ;
      VIA 31.038 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.033 31.083 31.067 ;
      VIA 31.038 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 30.493 31.083 30.527 ;
      VIA 31.038 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.953 31.083 29.987 ;
      VIA 31.038 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.413 31.083 29.447 ;
      VIA 31.038 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.873 31.083 28.907 ;
      VIA 31.038 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.333 31.083 28.367 ;
      VIA 31.038 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.793 31.083 27.827 ;
      VIA 31.038 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.253 31.083 27.287 ;
      VIA 31.038 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.713 31.083 26.747 ;
      VIA 31.038 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.173 31.083 26.207 ;
      VIA 31.038 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.633 31.083 25.667 ;
      VIA 31.038 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.093 31.083 25.127 ;
      VIA 31.038 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.553 31.083 24.587 ;
      VIA 31.038 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.013 31.083 24.047 ;
      VIA 31.038 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 23.473 31.083 23.507 ;
      VIA 31.038 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.933 31.083 22.967 ;
      VIA 31.038 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.393 31.083 22.427 ;
      VIA 31.038 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.853 31.083 21.887 ;
      VIA 31.038 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.313 31.083 21.347 ;
      VIA 31.038 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.773 31.083 20.807 ;
      VIA 31.038 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.233 31.083 20.267 ;
      VIA 31.038 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.693 31.083 19.727 ;
      VIA 31.038 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.153 31.083 19.187 ;
      VIA 31.038 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.613 31.083 18.647 ;
      VIA 31.038 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.073 31.083 18.107 ;
      VIA 31.038 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 17.533 31.083 17.567 ;
      VIA 31.038 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.993 31.083 17.027 ;
      VIA 31.038 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.453 31.083 16.487 ;
      VIA 31.038 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.913 31.083 15.947 ;
      VIA 31.038 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.373 31.083 15.407 ;
      VIA 31.038 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.833 31.083 14.867 ;
      VIA 31.038 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.293 31.083 14.327 ;
      VIA 31.038 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.753 31.083 13.787 ;
      VIA 31.038 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.213 31.083 13.247 ;
      VIA 31.038 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.673 31.083 12.707 ;
      VIA 31.038 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.133 31.083 12.167 ;
      VIA 31.038 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.593 31.083 11.627 ;
      VIA 31.038 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.053 31.083 11.087 ;
      VIA 31.038 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 10.513 31.083 10.547 ;
      VIA 31.038 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.973 31.083 10.007 ;
      VIA 31.038 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.433 31.083 9.467 ;
      VIA 31.038 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.893 31.083 8.927 ;
      VIA 31.038 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.353 31.083 8.387 ;
      VIA 31.038 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.813 31.083 7.847 ;
      VIA 31.038 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.273 31.083 7.307 ;
      VIA 31.038 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.733 31.083 6.767 ;
      VIA 31.038 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.193 31.083 6.227 ;
      VIA 31.038 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.653 31.083 5.687 ;
      VIA 31.038 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.113 31.083 5.147 ;
      VIA 31.038 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.573 31.083 4.607 ;
      VIA 31.038 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.033 31.083 4.067 ;
      VIA 31.038 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 3.493 31.083 3.527 ;
      VIA 31.038 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.953 31.083 2.987 ;
      VIA 31.038 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.413 31.083 2.447 ;
      VIA 31.038 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.873 31.083 1.907 ;
      VIA 31.038 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.333 31.083 1.367 ;
      VIA 31.038 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 58.033 25.179 58.067 ;
      VIA 25.134 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 57.493 25.179 57.527 ;
      VIA 25.134 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 56.953 25.179 56.987 ;
      VIA 25.134 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 56.413 25.179 56.447 ;
      VIA 25.134 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 55.873 25.179 55.907 ;
      VIA 25.134 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 55.333 25.179 55.367 ;
      VIA 25.134 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 54.793 25.179 54.827 ;
      VIA 25.134 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 54.253 25.179 54.287 ;
      VIA 25.134 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 53.713 25.179 53.747 ;
      VIA 25.134 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 53.173 25.179 53.207 ;
      VIA 25.134 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 52.633 25.179 52.667 ;
      VIA 25.134 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 52.093 25.179 52.127 ;
      VIA 25.134 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 51.553 25.179 51.587 ;
      VIA 25.134 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 51.013 25.179 51.047 ;
      VIA 25.134 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 50.473 25.179 50.507 ;
      VIA 25.134 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 49.933 25.179 49.967 ;
      VIA 25.134 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 49.393 25.179 49.427 ;
      VIA 25.134 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 48.853 25.179 48.887 ;
      VIA 25.134 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 48.313 25.179 48.347 ;
      VIA 25.134 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 47.773 25.179 47.807 ;
      VIA 25.134 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 47.233 25.179 47.267 ;
      VIA 25.134 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 46.693 25.179 46.727 ;
      VIA 25.134 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 46.153 25.179 46.187 ;
      VIA 25.134 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 45.613 25.179 45.647 ;
      VIA 25.134 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 45.073 25.179 45.107 ;
      VIA 25.134 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 44.533 25.179 44.567 ;
      VIA 25.134 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 43.993 25.179 44.027 ;
      VIA 25.134 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 43.453 25.179 43.487 ;
      VIA 25.134 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 42.913 25.179 42.947 ;
      VIA 25.134 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 42.373 25.179 42.407 ;
      VIA 25.134 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 41.833 25.179 41.867 ;
      VIA 25.134 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 41.293 25.179 41.327 ;
      VIA 25.134 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 40.753 25.179 40.787 ;
      VIA 25.134 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 40.213 25.179 40.247 ;
      VIA 25.134 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.673 25.179 39.707 ;
      VIA 25.134 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.133 25.179 39.167 ;
      VIA 25.134 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.593 25.179 38.627 ;
      VIA 25.134 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.053 25.179 38.087 ;
      VIA 25.134 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 37.513 25.179 37.547 ;
      VIA 25.134 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.973 25.179 37.007 ;
      VIA 25.134 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.433 25.179 36.467 ;
      VIA 25.134 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.893 25.179 35.927 ;
      VIA 25.134 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.353 25.179 35.387 ;
      VIA 25.134 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.813 25.179 34.847 ;
      VIA 25.134 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.273 25.179 34.307 ;
      VIA 25.134 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.733 25.179 33.767 ;
      VIA 25.134 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.193 25.179 33.227 ;
      VIA 25.134 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.653 25.179 32.687 ;
      VIA 25.134 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.113 25.179 32.147 ;
      VIA 25.134 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.573 25.179 31.607 ;
      VIA 25.134 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.033 25.179 31.067 ;
      VIA 25.134 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 30.493 25.179 30.527 ;
      VIA 25.134 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.953 25.179 29.987 ;
      VIA 25.134 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.413 25.179 29.447 ;
      VIA 25.134 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.873 25.179 28.907 ;
      VIA 25.134 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.333 25.179 28.367 ;
      VIA 25.134 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.793 25.179 27.827 ;
      VIA 25.134 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.253 25.179 27.287 ;
      VIA 25.134 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.713 25.179 26.747 ;
      VIA 25.134 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.173 25.179 26.207 ;
      VIA 25.134 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.633 25.179 25.667 ;
      VIA 25.134 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.093 25.179 25.127 ;
      VIA 25.134 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.553 25.179 24.587 ;
      VIA 25.134 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.013 25.179 24.047 ;
      VIA 25.134 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 23.473 25.179 23.507 ;
      VIA 25.134 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.933 25.179 22.967 ;
      VIA 25.134 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.393 25.179 22.427 ;
      VIA 25.134 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.853 25.179 21.887 ;
      VIA 25.134 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.313 25.179 21.347 ;
      VIA 25.134 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.773 25.179 20.807 ;
      VIA 25.134 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.233 25.179 20.267 ;
      VIA 25.134 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.693 25.179 19.727 ;
      VIA 25.134 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.153 25.179 19.187 ;
      VIA 25.134 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.613 25.179 18.647 ;
      VIA 25.134 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.073 25.179 18.107 ;
      VIA 25.134 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 17.533 25.179 17.567 ;
      VIA 25.134 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.993 25.179 17.027 ;
      VIA 25.134 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.453 25.179 16.487 ;
      VIA 25.134 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.913 25.179 15.947 ;
      VIA 25.134 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.373 25.179 15.407 ;
      VIA 25.134 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.833 25.179 14.867 ;
      VIA 25.134 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.293 25.179 14.327 ;
      VIA 25.134 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.753 25.179 13.787 ;
      VIA 25.134 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.213 25.179 13.247 ;
      VIA 25.134 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.673 25.179 12.707 ;
      VIA 25.134 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.133 25.179 12.167 ;
      VIA 25.134 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.593 25.179 11.627 ;
      VIA 25.134 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.053 25.179 11.087 ;
      VIA 25.134 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 10.513 25.179 10.547 ;
      VIA 25.134 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.973 25.179 10.007 ;
      VIA 25.134 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.433 25.179 9.467 ;
      VIA 25.134 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.893 25.179 8.927 ;
      VIA 25.134 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.353 25.179 8.387 ;
      VIA 25.134 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.813 25.179 7.847 ;
      VIA 25.134 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.273 25.179 7.307 ;
      VIA 25.134 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.733 25.179 6.767 ;
      VIA 25.134 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.193 25.179 6.227 ;
      VIA 25.134 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.653 25.179 5.687 ;
      VIA 25.134 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.113 25.179 5.147 ;
      VIA 25.134 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.573 25.179 4.607 ;
      VIA 25.134 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.033 25.179 4.067 ;
      VIA 25.134 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 3.493 25.179 3.527 ;
      VIA 25.134 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.953 25.179 2.987 ;
      VIA 25.134 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.413 25.179 2.447 ;
      VIA 25.134 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.873 25.179 1.907 ;
      VIA 25.134 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.333 25.179 1.367 ;
      VIA 25.134 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 58.033 19.275 58.067 ;
      VIA 19.23 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 57.493 19.275 57.527 ;
      VIA 19.23 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 56.953 19.275 56.987 ;
      VIA 19.23 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 56.413 19.275 56.447 ;
      VIA 19.23 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 55.873 19.275 55.907 ;
      VIA 19.23 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 55.333 19.275 55.367 ;
      VIA 19.23 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 54.793 19.275 54.827 ;
      VIA 19.23 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 54.253 19.275 54.287 ;
      VIA 19.23 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 53.713 19.275 53.747 ;
      VIA 19.23 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 53.173 19.275 53.207 ;
      VIA 19.23 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 52.633 19.275 52.667 ;
      VIA 19.23 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 52.093 19.275 52.127 ;
      VIA 19.23 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 51.553 19.275 51.587 ;
      VIA 19.23 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 51.013 19.275 51.047 ;
      VIA 19.23 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 50.473 19.275 50.507 ;
      VIA 19.23 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 49.933 19.275 49.967 ;
      VIA 19.23 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 49.393 19.275 49.427 ;
      VIA 19.23 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 48.853 19.275 48.887 ;
      VIA 19.23 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 48.313 19.275 48.347 ;
      VIA 19.23 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 47.773 19.275 47.807 ;
      VIA 19.23 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 47.233 19.275 47.267 ;
      VIA 19.23 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 46.693 19.275 46.727 ;
      VIA 19.23 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 46.153 19.275 46.187 ;
      VIA 19.23 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 45.613 19.275 45.647 ;
      VIA 19.23 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 45.073 19.275 45.107 ;
      VIA 19.23 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 44.533 19.275 44.567 ;
      VIA 19.23 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 43.993 19.275 44.027 ;
      VIA 19.23 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 43.453 19.275 43.487 ;
      VIA 19.23 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 42.913 19.275 42.947 ;
      VIA 19.23 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 42.373 19.275 42.407 ;
      VIA 19.23 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 41.833 19.275 41.867 ;
      VIA 19.23 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 41.293 19.275 41.327 ;
      VIA 19.23 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 40.753 19.275 40.787 ;
      VIA 19.23 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 40.213 19.275 40.247 ;
      VIA 19.23 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.673 19.275 39.707 ;
      VIA 19.23 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.133 19.275 39.167 ;
      VIA 19.23 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.593 19.275 38.627 ;
      VIA 19.23 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.053 19.275 38.087 ;
      VIA 19.23 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 37.513 19.275 37.547 ;
      VIA 19.23 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.973 19.275 37.007 ;
      VIA 19.23 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.433 19.275 36.467 ;
      VIA 19.23 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.893 19.275 35.927 ;
      VIA 19.23 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.353 19.275 35.387 ;
      VIA 19.23 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.813 19.275 34.847 ;
      VIA 19.23 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.273 19.275 34.307 ;
      VIA 19.23 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.733 19.275 33.767 ;
      VIA 19.23 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.193 19.275 33.227 ;
      VIA 19.23 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.653 19.275 32.687 ;
      VIA 19.23 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.113 19.275 32.147 ;
      VIA 19.23 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.573 19.275 31.607 ;
      VIA 19.23 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.033 19.275 31.067 ;
      VIA 19.23 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 30.493 19.275 30.527 ;
      VIA 19.23 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.953 19.275 29.987 ;
      VIA 19.23 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.413 19.275 29.447 ;
      VIA 19.23 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.873 19.275 28.907 ;
      VIA 19.23 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.333 19.275 28.367 ;
      VIA 19.23 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.793 19.275 27.827 ;
      VIA 19.23 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.253 19.275 27.287 ;
      VIA 19.23 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.713 19.275 26.747 ;
      VIA 19.23 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.173 19.275 26.207 ;
      VIA 19.23 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.633 19.275 25.667 ;
      VIA 19.23 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.093 19.275 25.127 ;
      VIA 19.23 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.553 19.275 24.587 ;
      VIA 19.23 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.013 19.275 24.047 ;
      VIA 19.23 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 23.473 19.275 23.507 ;
      VIA 19.23 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.933 19.275 22.967 ;
      VIA 19.23 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.393 19.275 22.427 ;
      VIA 19.23 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.853 19.275 21.887 ;
      VIA 19.23 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.313 19.275 21.347 ;
      VIA 19.23 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.773 19.275 20.807 ;
      VIA 19.23 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.233 19.275 20.267 ;
      VIA 19.23 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.693 19.275 19.727 ;
      VIA 19.23 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.153 19.275 19.187 ;
      VIA 19.23 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.613 19.275 18.647 ;
      VIA 19.23 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.073 19.275 18.107 ;
      VIA 19.23 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 17.533 19.275 17.567 ;
      VIA 19.23 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.993 19.275 17.027 ;
      VIA 19.23 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.453 19.275 16.487 ;
      VIA 19.23 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.913 19.275 15.947 ;
      VIA 19.23 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.373 19.275 15.407 ;
      VIA 19.23 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.833 19.275 14.867 ;
      VIA 19.23 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.293 19.275 14.327 ;
      VIA 19.23 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.753 19.275 13.787 ;
      VIA 19.23 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.213 19.275 13.247 ;
      VIA 19.23 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.673 19.275 12.707 ;
      VIA 19.23 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.133 19.275 12.167 ;
      VIA 19.23 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.593 19.275 11.627 ;
      VIA 19.23 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.053 19.275 11.087 ;
      VIA 19.23 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 10.513 19.275 10.547 ;
      VIA 19.23 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.973 19.275 10.007 ;
      VIA 19.23 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.433 19.275 9.467 ;
      VIA 19.23 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.893 19.275 8.927 ;
      VIA 19.23 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.353 19.275 8.387 ;
      VIA 19.23 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.813 19.275 7.847 ;
      VIA 19.23 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.273 19.275 7.307 ;
      VIA 19.23 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.733 19.275 6.767 ;
      VIA 19.23 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.193 19.275 6.227 ;
      VIA 19.23 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.653 19.275 5.687 ;
      VIA 19.23 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.113 19.275 5.147 ;
      VIA 19.23 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.573 19.275 4.607 ;
      VIA 19.23 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.033 19.275 4.067 ;
      VIA 19.23 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 3.493 19.275 3.527 ;
      VIA 19.23 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.953 19.275 2.987 ;
      VIA 19.23 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.413 19.275 2.447 ;
      VIA 19.23 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.873 19.275 1.907 ;
      VIA 19.23 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.333 19.275 1.367 ;
      VIA 19.23 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 58.033 13.371 58.067 ;
      VIA 13.326 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 57.493 13.371 57.527 ;
      VIA 13.326 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 56.953 13.371 56.987 ;
      VIA 13.326 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 56.413 13.371 56.447 ;
      VIA 13.326 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 55.873 13.371 55.907 ;
      VIA 13.326 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 55.333 13.371 55.367 ;
      VIA 13.326 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 54.793 13.371 54.827 ;
      VIA 13.326 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 54.253 13.371 54.287 ;
      VIA 13.326 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 53.713 13.371 53.747 ;
      VIA 13.326 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 53.173 13.371 53.207 ;
      VIA 13.326 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 52.633 13.371 52.667 ;
      VIA 13.326 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 52.093 13.371 52.127 ;
      VIA 13.326 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 51.553 13.371 51.587 ;
      VIA 13.326 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 51.013 13.371 51.047 ;
      VIA 13.326 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 50.473 13.371 50.507 ;
      VIA 13.326 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 49.933 13.371 49.967 ;
      VIA 13.326 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 49.393 13.371 49.427 ;
      VIA 13.326 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 48.853 13.371 48.887 ;
      VIA 13.326 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 48.313 13.371 48.347 ;
      VIA 13.326 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 47.773 13.371 47.807 ;
      VIA 13.326 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 47.233 13.371 47.267 ;
      VIA 13.326 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 46.693 13.371 46.727 ;
      VIA 13.326 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 46.153 13.371 46.187 ;
      VIA 13.326 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 45.613 13.371 45.647 ;
      VIA 13.326 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 45.073 13.371 45.107 ;
      VIA 13.326 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 44.533 13.371 44.567 ;
      VIA 13.326 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 43.993 13.371 44.027 ;
      VIA 13.326 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 43.453 13.371 43.487 ;
      VIA 13.326 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 42.913 13.371 42.947 ;
      VIA 13.326 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 42.373 13.371 42.407 ;
      VIA 13.326 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 41.833 13.371 41.867 ;
      VIA 13.326 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 41.293 13.371 41.327 ;
      VIA 13.326 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 40.753 13.371 40.787 ;
      VIA 13.326 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 40.213 13.371 40.247 ;
      VIA 13.326 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.673 13.371 39.707 ;
      VIA 13.326 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.133 13.371 39.167 ;
      VIA 13.326 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.593 13.371 38.627 ;
      VIA 13.326 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.053 13.371 38.087 ;
      VIA 13.326 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 37.513 13.371 37.547 ;
      VIA 13.326 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.973 13.371 37.007 ;
      VIA 13.326 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.433 13.371 36.467 ;
      VIA 13.326 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.893 13.371 35.927 ;
      VIA 13.326 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.353 13.371 35.387 ;
      VIA 13.326 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.813 13.371 34.847 ;
      VIA 13.326 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.273 13.371 34.307 ;
      VIA 13.326 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.733 13.371 33.767 ;
      VIA 13.326 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.193 13.371 33.227 ;
      VIA 13.326 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.653 13.371 32.687 ;
      VIA 13.326 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.113 13.371 32.147 ;
      VIA 13.326 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.573 13.371 31.607 ;
      VIA 13.326 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.033 13.371 31.067 ;
      VIA 13.326 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 30.493 13.371 30.527 ;
      VIA 13.326 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.953 13.371 29.987 ;
      VIA 13.326 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.413 13.371 29.447 ;
      VIA 13.326 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.873 13.371 28.907 ;
      VIA 13.326 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.333 13.371 28.367 ;
      VIA 13.326 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.793 13.371 27.827 ;
      VIA 13.326 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.253 13.371 27.287 ;
      VIA 13.326 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.713 13.371 26.747 ;
      VIA 13.326 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.173 13.371 26.207 ;
      VIA 13.326 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.633 13.371 25.667 ;
      VIA 13.326 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.093 13.371 25.127 ;
      VIA 13.326 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.553 13.371 24.587 ;
      VIA 13.326 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.013 13.371 24.047 ;
      VIA 13.326 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 23.473 13.371 23.507 ;
      VIA 13.326 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.933 13.371 22.967 ;
      VIA 13.326 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.393 13.371 22.427 ;
      VIA 13.326 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.853 13.371 21.887 ;
      VIA 13.326 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.313 13.371 21.347 ;
      VIA 13.326 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.773 13.371 20.807 ;
      VIA 13.326 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.233 13.371 20.267 ;
      VIA 13.326 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.693 13.371 19.727 ;
      VIA 13.326 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.153 13.371 19.187 ;
      VIA 13.326 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.613 13.371 18.647 ;
      VIA 13.326 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.073 13.371 18.107 ;
      VIA 13.326 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 17.533 13.371 17.567 ;
      VIA 13.326 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.993 13.371 17.027 ;
      VIA 13.326 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.453 13.371 16.487 ;
      VIA 13.326 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.913 13.371 15.947 ;
      VIA 13.326 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.373 13.371 15.407 ;
      VIA 13.326 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.833 13.371 14.867 ;
      VIA 13.326 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.293 13.371 14.327 ;
      VIA 13.326 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.753 13.371 13.787 ;
      VIA 13.326 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.213 13.371 13.247 ;
      VIA 13.326 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.673 13.371 12.707 ;
      VIA 13.326 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.133 13.371 12.167 ;
      VIA 13.326 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.593 13.371 11.627 ;
      VIA 13.326 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.053 13.371 11.087 ;
      VIA 13.326 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 10.513 13.371 10.547 ;
      VIA 13.326 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.973 13.371 10.007 ;
      VIA 13.326 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.433 13.371 9.467 ;
      VIA 13.326 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.893 13.371 8.927 ;
      VIA 13.326 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.353 13.371 8.387 ;
      VIA 13.326 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.813 13.371 7.847 ;
      VIA 13.326 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.273 13.371 7.307 ;
      VIA 13.326 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.733 13.371 6.767 ;
      VIA 13.326 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.193 13.371 6.227 ;
      VIA 13.326 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.653 13.371 5.687 ;
      VIA 13.326 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.113 13.371 5.147 ;
      VIA 13.326 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.573 13.371 4.607 ;
      VIA 13.326 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.033 13.371 4.067 ;
      VIA 13.326 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 3.493 13.371 3.527 ;
      VIA 13.326 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.953 13.371 2.987 ;
      VIA 13.326 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.413 13.371 2.447 ;
      VIA 13.326 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.873 13.371 1.907 ;
      VIA 13.326 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.333 13.371 1.367 ;
      VIA 13.326 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 58.033 7.467 58.067 ;
      VIA 7.422 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 57.493 7.467 57.527 ;
      VIA 7.422 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 56.953 7.467 56.987 ;
      VIA 7.422 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 56.413 7.467 56.447 ;
      VIA 7.422 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 55.873 7.467 55.907 ;
      VIA 7.422 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 55.333 7.467 55.367 ;
      VIA 7.422 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 54.793 7.467 54.827 ;
      VIA 7.422 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 54.253 7.467 54.287 ;
      VIA 7.422 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 53.713 7.467 53.747 ;
      VIA 7.422 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 53.173 7.467 53.207 ;
      VIA 7.422 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 52.633 7.467 52.667 ;
      VIA 7.422 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 52.093 7.467 52.127 ;
      VIA 7.422 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 51.553 7.467 51.587 ;
      VIA 7.422 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 51.013 7.467 51.047 ;
      VIA 7.422 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 50.473 7.467 50.507 ;
      VIA 7.422 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 49.933 7.467 49.967 ;
      VIA 7.422 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 49.393 7.467 49.427 ;
      VIA 7.422 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 48.853 7.467 48.887 ;
      VIA 7.422 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 48.313 7.467 48.347 ;
      VIA 7.422 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 47.773 7.467 47.807 ;
      VIA 7.422 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 47.233 7.467 47.267 ;
      VIA 7.422 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 46.693 7.467 46.727 ;
      VIA 7.422 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 46.153 7.467 46.187 ;
      VIA 7.422 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 45.613 7.467 45.647 ;
      VIA 7.422 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 45.073 7.467 45.107 ;
      VIA 7.422 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 44.533 7.467 44.567 ;
      VIA 7.422 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 43.993 7.467 44.027 ;
      VIA 7.422 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 43.453 7.467 43.487 ;
      VIA 7.422 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 42.913 7.467 42.947 ;
      VIA 7.422 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 42.373 7.467 42.407 ;
      VIA 7.422 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 41.833 7.467 41.867 ;
      VIA 7.422 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 41.293 7.467 41.327 ;
      VIA 7.422 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 40.753 7.467 40.787 ;
      VIA 7.422 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 40.213 7.467 40.247 ;
      VIA 7.422 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.673 7.467 39.707 ;
      VIA 7.422 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.133 7.467 39.167 ;
      VIA 7.422 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.593 7.467 38.627 ;
      VIA 7.422 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.053 7.467 38.087 ;
      VIA 7.422 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 37.513 7.467 37.547 ;
      VIA 7.422 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.973 7.467 37.007 ;
      VIA 7.422 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.433 7.467 36.467 ;
      VIA 7.422 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.893 7.467 35.927 ;
      VIA 7.422 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.353 7.467 35.387 ;
      VIA 7.422 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.813 7.467 34.847 ;
      VIA 7.422 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.273 7.467 34.307 ;
      VIA 7.422 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.733 7.467 33.767 ;
      VIA 7.422 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.193 7.467 33.227 ;
      VIA 7.422 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.653 7.467 32.687 ;
      VIA 7.422 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.113 7.467 32.147 ;
      VIA 7.422 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.573 7.467 31.607 ;
      VIA 7.422 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.033 7.467 31.067 ;
      VIA 7.422 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 30.493 7.467 30.527 ;
      VIA 7.422 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.953 7.467 29.987 ;
      VIA 7.422 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.413 7.467 29.447 ;
      VIA 7.422 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.873 7.467 28.907 ;
      VIA 7.422 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.333 7.467 28.367 ;
      VIA 7.422 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.793 7.467 27.827 ;
      VIA 7.422 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.253 7.467 27.287 ;
      VIA 7.422 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.713 7.467 26.747 ;
      VIA 7.422 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.173 7.467 26.207 ;
      VIA 7.422 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.633 7.467 25.667 ;
      VIA 7.422 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.093 7.467 25.127 ;
      VIA 7.422 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.553 7.467 24.587 ;
      VIA 7.422 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.013 7.467 24.047 ;
      VIA 7.422 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 23.473 7.467 23.507 ;
      VIA 7.422 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.933 7.467 22.967 ;
      VIA 7.422 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.393 7.467 22.427 ;
      VIA 7.422 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.853 7.467 21.887 ;
      VIA 7.422 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.313 7.467 21.347 ;
      VIA 7.422 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.773 7.467 20.807 ;
      VIA 7.422 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.233 7.467 20.267 ;
      VIA 7.422 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.693 7.467 19.727 ;
      VIA 7.422 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.153 7.467 19.187 ;
      VIA 7.422 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.613 7.467 18.647 ;
      VIA 7.422 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.073 7.467 18.107 ;
      VIA 7.422 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 17.533 7.467 17.567 ;
      VIA 7.422 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.993 7.467 17.027 ;
      VIA 7.422 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.453 7.467 16.487 ;
      VIA 7.422 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.913 7.467 15.947 ;
      VIA 7.422 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.373 7.467 15.407 ;
      VIA 7.422 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.833 7.467 14.867 ;
      VIA 7.422 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.293 7.467 14.327 ;
      VIA 7.422 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.753 7.467 13.787 ;
      VIA 7.422 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.213 7.467 13.247 ;
      VIA 7.422 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.673 7.467 12.707 ;
      VIA 7.422 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.133 7.467 12.167 ;
      VIA 7.422 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.593 7.467 11.627 ;
      VIA 7.422 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.053 7.467 11.087 ;
      VIA 7.422 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 10.513 7.467 10.547 ;
      VIA 7.422 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.973 7.467 10.007 ;
      VIA 7.422 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.433 7.467 9.467 ;
      VIA 7.422 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.893 7.467 8.927 ;
      VIA 7.422 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.353 7.467 8.387 ;
      VIA 7.422 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.813 7.467 7.847 ;
      VIA 7.422 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.273 7.467 7.307 ;
      VIA 7.422 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.733 7.467 6.767 ;
      VIA 7.422 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.193 7.467 6.227 ;
      VIA 7.422 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.653 7.467 5.687 ;
      VIA 7.422 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.113 7.467 5.147 ;
      VIA 7.422 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.573 7.467 4.607 ;
      VIA 7.422 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.033 7.467 4.067 ;
      VIA 7.422 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 3.493 7.467 3.527 ;
      VIA 7.422 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.953 7.467 2.987 ;
      VIA 7.422 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.413 7.467 2.447 ;
      VIA 7.422 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.873 7.467 1.907 ;
      VIA 7.422 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.333 7.467 1.367 ;
      VIA 7.422 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 58.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 58.033 1.563 58.067 ;
      VIA 1.518 58.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 58.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 57.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 57.493 1.563 57.527 ;
      VIA 1.518 57.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 57.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 56.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 56.953 1.563 56.987 ;
      VIA 1.518 56.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 56.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 56.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 56.413 1.563 56.447 ;
      VIA 1.518 56.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 56.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 55.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 55.873 1.563 55.907 ;
      VIA 1.518 55.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 55.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 55.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 55.333 1.563 55.367 ;
      VIA 1.518 55.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 55.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 54.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 54.793 1.563 54.827 ;
      VIA 1.518 54.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 54.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 54.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 54.253 1.563 54.287 ;
      VIA 1.518 54.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 54.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 53.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 53.713 1.563 53.747 ;
      VIA 1.518 53.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 53.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 53.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 53.173 1.563 53.207 ;
      VIA 1.518 53.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 53.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 52.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 52.633 1.563 52.667 ;
      VIA 1.518 52.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 52.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 52.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 52.093 1.563 52.127 ;
      VIA 1.518 52.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 52.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 51.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 51.553 1.563 51.587 ;
      VIA 1.518 51.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 51.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 51.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 51.013 1.563 51.047 ;
      VIA 1.518 51.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 51.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 50.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 50.473 1.563 50.507 ;
      VIA 1.518 50.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 50.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 49.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 49.933 1.563 49.967 ;
      VIA 1.518 49.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 49.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 49.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 49.393 1.563 49.427 ;
      VIA 1.518 49.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 49.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 48.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 48.853 1.563 48.887 ;
      VIA 1.518 48.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 48.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 48.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 48.313 1.563 48.347 ;
      VIA 1.518 48.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 48.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 47.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 47.773 1.563 47.807 ;
      VIA 1.518 47.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 47.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 47.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 47.233 1.563 47.267 ;
      VIA 1.518 47.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 47.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 46.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 46.693 1.563 46.727 ;
      VIA 1.518 46.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 46.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 46.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 46.153 1.563 46.187 ;
      VIA 1.518 46.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 46.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 45.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 45.613 1.563 45.647 ;
      VIA 1.518 45.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 45.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 45.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 45.073 1.563 45.107 ;
      VIA 1.518 45.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 45.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 44.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 44.533 1.563 44.567 ;
      VIA 1.518 44.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 44.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 44.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 43.993 1.563 44.027 ;
      VIA 1.518 44.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 44.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 43.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 43.453 1.563 43.487 ;
      VIA 1.518 43.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 43.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 42.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 42.913 1.563 42.947 ;
      VIA 1.518 42.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 42.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 42.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 42.373 1.563 42.407 ;
      VIA 1.518 42.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 42.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 41.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 41.833 1.563 41.867 ;
      VIA 1.518 41.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 41.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 41.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 41.293 1.563 41.327 ;
      VIA 1.518 41.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 41.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 40.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 40.753 1.563 40.787 ;
      VIA 1.518 40.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 40.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 40.213 1.563 40.247 ;
      VIA 1.518 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.673 1.563 39.707 ;
      VIA 1.518 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.133 1.563 39.167 ;
      VIA 1.518 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.593 1.563 38.627 ;
      VIA 1.518 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.053 1.563 38.087 ;
      VIA 1.518 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 37.513 1.563 37.547 ;
      VIA 1.518 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.973 1.563 37.007 ;
      VIA 1.518 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.433 1.563 36.467 ;
      VIA 1.518 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.893 1.563 35.927 ;
      VIA 1.518 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.353 1.563 35.387 ;
      VIA 1.518 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.813 1.563 34.847 ;
      VIA 1.518 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.273 1.563 34.307 ;
      VIA 1.518 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.733 1.563 33.767 ;
      VIA 1.518 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.193 1.563 33.227 ;
      VIA 1.518 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.653 1.563 32.687 ;
      VIA 1.518 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.113 1.563 32.147 ;
      VIA 1.518 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.573 1.563 31.607 ;
      VIA 1.518 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.033 1.563 31.067 ;
      VIA 1.518 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 30.493 1.563 30.527 ;
      VIA 1.518 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.953 1.563 29.987 ;
      VIA 1.518 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.413 1.563 29.447 ;
      VIA 1.518 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.873 1.563 28.907 ;
      VIA 1.518 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.333 1.563 28.367 ;
      VIA 1.518 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.793 1.563 27.827 ;
      VIA 1.518 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.253 1.563 27.287 ;
      VIA 1.518 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.713 1.563 26.747 ;
      VIA 1.518 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.173 1.563 26.207 ;
      VIA 1.518 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.633 1.563 25.667 ;
      VIA 1.518 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.093 1.563 25.127 ;
      VIA 1.518 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.553 1.563 24.587 ;
      VIA 1.518 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.013 1.563 24.047 ;
      VIA 1.518 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 23.473 1.563 23.507 ;
      VIA 1.518 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.933 1.563 22.967 ;
      VIA 1.518 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.393 1.563 22.427 ;
      VIA 1.518 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.853 1.563 21.887 ;
      VIA 1.518 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.313 1.563 21.347 ;
      VIA 1.518 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.773 1.563 20.807 ;
      VIA 1.518 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.233 1.563 20.267 ;
      VIA 1.518 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.693 1.563 19.727 ;
      VIA 1.518 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.153 1.563 19.187 ;
      VIA 1.518 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.613 1.563 18.647 ;
      VIA 1.518 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.073 1.563 18.107 ;
      VIA 1.518 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 17.533 1.563 17.567 ;
      VIA 1.518 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.993 1.563 17.027 ;
      VIA 1.518 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.453 1.563 16.487 ;
      VIA 1.518 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.913 1.563 15.947 ;
      VIA 1.518 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.373 1.563 15.407 ;
      VIA 1.518 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.833 1.563 14.867 ;
      VIA 1.518 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.293 1.563 14.327 ;
      VIA 1.518 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.753 1.563 13.787 ;
      VIA 1.518 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.213 1.563 13.247 ;
      VIA 1.518 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.673 1.563 12.707 ;
      VIA 1.518 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.133 1.563 12.167 ;
      VIA 1.518 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.593 1.563 11.627 ;
      VIA 1.518 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.053 1.563 11.087 ;
      VIA 1.518 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 10.513 1.563 10.547 ;
      VIA 1.518 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.973 1.563 10.007 ;
      VIA 1.518 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.433 1.563 9.467 ;
      VIA 1.518 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.893 1.563 8.927 ;
      VIA 1.518 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.353 1.563 8.387 ;
      VIA 1.518 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.813 1.563 7.847 ;
      VIA 1.518 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.273 1.563 7.307 ;
      VIA 1.518 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.733 1.563 6.767 ;
      VIA 1.518 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.193 1.563 6.227 ;
      VIA 1.518 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.653 1.563 5.687 ;
      VIA 1.518 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.113 1.563 5.147 ;
      VIA 1.518 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 29.565 58.05 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 57.51 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 56.97 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 56.43 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 55.89 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 55.35 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 54.81 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 54.27 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 53.73 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 53.19 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 52.65 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 52.11 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 51.57 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 51.03 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 50.49 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 49.95 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 49.41 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 48.87 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 48.33 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 47.79 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 47.25 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 46.71 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 46.17 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 45.63 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 45.09 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 44.55 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 44.01 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 43.47 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 42.93 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 42.39 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 41.85 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 41.31 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 40.77 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 40.23 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 39.69 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 39.15 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 38.61 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 38.07 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 37.53 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 36.99 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 36.45 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 35.91 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 35.37 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 34.83 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 34.29 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 33.75 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 33.21 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 32.67 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 32.13 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 31.59 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 31.05 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 30.51 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 29.97 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 29.43 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 28.89 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 28.35 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 27.81 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 27.27 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 26.73 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 26.19 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 25.65 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 25.11 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 24.57 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 24.03 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 23.49 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 22.95 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 22.41 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 21.87 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 21.33 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 20.79 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 20.25 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 19.71 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 19.17 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 18.63 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 18.09 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 17.55 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 17.01 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 16.47 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 15.93 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 15.39 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 14.85 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 14.31 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 13.77 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 13.23 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 12.69 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 12.15 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 11.61 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 11.07 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 10.53 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 9.99 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 9.45 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 8.91 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 8.37 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 7.83 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 7.29 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 6.75 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 6.21 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 5.67 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 5.13 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 4.59 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 4.05 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 3.51 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 2.97 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 2.43 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 1.89 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 1.35 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.266 55.449 54.522 55.737 ;
        RECT  1.266 49.449 54.522 49.737 ;
        RECT  1.266 43.449 54.522 43.737 ;
        RECT  1.266 37.449 54.522 37.737 ;
        RECT  1.266 31.449 54.522 31.737 ;
        RECT  1.266 25.449 54.522 25.737 ;
        RECT  1.266 19.449 54.522 19.737 ;
        RECT  1.266 13.449 54.522 13.737 ;
        RECT  1.266 7.449 54.522 7.737 ;
        RECT  1.266 1.449 54.522 1.737 ;
      LAYER M5 ;
        RECT  54.402 1.057 54.522 57.803 ;
        RECT  48.498 1.057 48.618 57.803 ;
        RECT  42.594 1.057 42.714 57.803 ;
        RECT  36.69 1.057 36.81 57.803 ;
        RECT  30.786 1.057 30.906 57.803 ;
        RECT  24.882 1.057 25.002 57.803 ;
        RECT  18.978 1.057 19.098 57.803 ;
        RECT  13.074 1.057 13.194 57.803 ;
        RECT  7.17 1.057 7.29 57.803 ;
        RECT  1.266 1.057 1.386 57.803 ;
      LAYER M2 ;
        RECT  1.026 57.771 58.104 57.789 ;
        RECT  1.026 57.231 58.104 57.249 ;
        RECT  1.026 56.691 58.104 56.709 ;
        RECT  1.026 56.151 58.104 56.169 ;
        RECT  1.026 55.611 58.104 55.629 ;
        RECT  1.026 55.071 58.104 55.089 ;
        RECT  1.026 54.531 58.104 54.549 ;
        RECT  1.026 53.991 58.104 54.009 ;
        RECT  1.026 53.451 58.104 53.469 ;
        RECT  1.026 52.911 58.104 52.929 ;
        RECT  1.026 52.371 58.104 52.389 ;
        RECT  1.026 51.831 58.104 51.849 ;
        RECT  1.026 51.291 58.104 51.309 ;
        RECT  1.026 50.751 58.104 50.769 ;
        RECT  1.026 50.211 58.104 50.229 ;
        RECT  1.026 49.671 58.104 49.689 ;
        RECT  1.026 49.131 58.104 49.149 ;
        RECT  1.026 48.591 58.104 48.609 ;
        RECT  1.026 48.051 58.104 48.069 ;
        RECT  1.026 47.511 58.104 47.529 ;
        RECT  1.026 46.971 58.104 46.989 ;
        RECT  1.026 46.431 58.104 46.449 ;
        RECT  1.026 45.891 58.104 45.909 ;
        RECT  1.026 45.351 58.104 45.369 ;
        RECT  1.026 44.811 58.104 44.829 ;
        RECT  1.026 44.271 58.104 44.289 ;
        RECT  1.026 43.731 58.104 43.749 ;
        RECT  1.026 43.191 58.104 43.209 ;
        RECT  1.026 42.651 58.104 42.669 ;
        RECT  1.026 42.111 58.104 42.129 ;
        RECT  1.026 41.571 58.104 41.589 ;
        RECT  1.026 41.031 58.104 41.049 ;
        RECT  1.026 40.491 58.104 40.509 ;
        RECT  1.026 39.951 58.104 39.969 ;
        RECT  1.026 39.411 58.104 39.429 ;
        RECT  1.026 38.871 58.104 38.889 ;
        RECT  1.026 38.331 58.104 38.349 ;
        RECT  1.026 37.791 58.104 37.809 ;
        RECT  1.026 37.251 58.104 37.269 ;
        RECT  1.026 36.711 58.104 36.729 ;
        RECT  1.026 36.171 58.104 36.189 ;
        RECT  1.026 35.631 58.104 35.649 ;
        RECT  1.026 35.091 58.104 35.109 ;
        RECT  1.026 34.551 58.104 34.569 ;
        RECT  1.026 34.011 58.104 34.029 ;
        RECT  1.026 33.471 58.104 33.489 ;
        RECT  1.026 32.931 58.104 32.949 ;
        RECT  1.026 32.391 58.104 32.409 ;
        RECT  1.026 31.851 58.104 31.869 ;
        RECT  1.026 31.311 58.104 31.329 ;
        RECT  1.026 30.771 58.104 30.789 ;
        RECT  1.026 30.231 58.104 30.249 ;
        RECT  1.026 29.691 58.104 29.709 ;
        RECT  1.026 29.151 58.104 29.169 ;
        RECT  1.026 28.611 58.104 28.629 ;
        RECT  1.026 28.071 58.104 28.089 ;
        RECT  1.026 27.531 58.104 27.549 ;
        RECT  1.026 26.991 58.104 27.009 ;
        RECT  1.026 26.451 58.104 26.469 ;
        RECT  1.026 25.911 58.104 25.929 ;
        RECT  1.026 25.371 58.104 25.389 ;
        RECT  1.026 24.831 58.104 24.849 ;
        RECT  1.026 24.291 58.104 24.309 ;
        RECT  1.026 23.751 58.104 23.769 ;
        RECT  1.026 23.211 58.104 23.229 ;
        RECT  1.026 22.671 58.104 22.689 ;
        RECT  1.026 22.131 58.104 22.149 ;
        RECT  1.026 21.591 58.104 21.609 ;
        RECT  1.026 21.051 58.104 21.069 ;
        RECT  1.026 20.511 58.104 20.529 ;
        RECT  1.026 19.971 58.104 19.989 ;
        RECT  1.026 19.431 58.104 19.449 ;
        RECT  1.026 18.891 58.104 18.909 ;
        RECT  1.026 18.351 58.104 18.369 ;
        RECT  1.026 17.811 58.104 17.829 ;
        RECT  1.026 17.271 58.104 17.289 ;
        RECT  1.026 16.731 58.104 16.749 ;
        RECT  1.026 16.191 58.104 16.209 ;
        RECT  1.026 15.651 58.104 15.669 ;
        RECT  1.026 15.111 58.104 15.129 ;
        RECT  1.026 14.571 58.104 14.589 ;
        RECT  1.026 14.031 58.104 14.049 ;
        RECT  1.026 13.491 58.104 13.509 ;
        RECT  1.026 12.951 58.104 12.969 ;
        RECT  1.026 12.411 58.104 12.429 ;
        RECT  1.026 11.871 58.104 11.889 ;
        RECT  1.026 11.331 58.104 11.349 ;
        RECT  1.026 10.791 58.104 10.809 ;
        RECT  1.026 10.251 58.104 10.269 ;
        RECT  1.026 9.711 58.104 9.729 ;
        RECT  1.026 9.171 58.104 9.189 ;
        RECT  1.026 8.631 58.104 8.649 ;
        RECT  1.026 8.091 58.104 8.109 ;
        RECT  1.026 7.551 58.104 7.569 ;
        RECT  1.026 7.011 58.104 7.029 ;
        RECT  1.026 6.471 58.104 6.489 ;
        RECT  1.026 5.931 58.104 5.949 ;
        RECT  1.026 5.391 58.104 5.409 ;
        RECT  1.026 4.851 58.104 4.869 ;
        RECT  1.026 4.311 58.104 4.329 ;
        RECT  1.026 3.771 58.104 3.789 ;
        RECT  1.026 3.231 58.104 3.249 ;
        RECT  1.026 2.691 58.104 2.709 ;
        RECT  1.026 2.151 58.104 2.169 ;
        RECT  1.026 1.611 58.104 1.629 ;
        RECT  1.026 1.071 58.104 1.089 ;
      LAYER M1 ;
        RECT  1.026 57.771 58.104 57.789 ;
        RECT  1.026 57.231 58.104 57.249 ;
        RECT  1.026 56.691 58.104 56.709 ;
        RECT  1.026 56.151 58.104 56.169 ;
        RECT  1.026 55.611 58.104 55.629 ;
        RECT  1.026 55.071 58.104 55.089 ;
        RECT  1.026 54.531 58.104 54.549 ;
        RECT  1.026 53.991 58.104 54.009 ;
        RECT  1.026 53.451 58.104 53.469 ;
        RECT  1.026 52.911 58.104 52.929 ;
        RECT  1.026 52.371 58.104 52.389 ;
        RECT  1.026 51.831 58.104 51.849 ;
        RECT  1.026 51.291 58.104 51.309 ;
        RECT  1.026 50.751 58.104 50.769 ;
        RECT  1.026 50.211 58.104 50.229 ;
        RECT  1.026 49.671 58.104 49.689 ;
        RECT  1.026 49.131 58.104 49.149 ;
        RECT  1.026 48.591 58.104 48.609 ;
        RECT  1.026 48.051 58.104 48.069 ;
        RECT  1.026 47.511 58.104 47.529 ;
        RECT  1.026 46.971 58.104 46.989 ;
        RECT  1.026 46.431 58.104 46.449 ;
        RECT  1.026 45.891 58.104 45.909 ;
        RECT  1.026 45.351 58.104 45.369 ;
        RECT  1.026 44.811 58.104 44.829 ;
        RECT  1.026 44.271 58.104 44.289 ;
        RECT  1.026 43.731 58.104 43.749 ;
        RECT  1.026 43.191 58.104 43.209 ;
        RECT  1.026 42.651 58.104 42.669 ;
        RECT  1.026 42.111 58.104 42.129 ;
        RECT  1.026 41.571 58.104 41.589 ;
        RECT  1.026 41.031 58.104 41.049 ;
        RECT  1.026 40.491 58.104 40.509 ;
        RECT  1.026 39.951 58.104 39.969 ;
        RECT  1.026 39.411 58.104 39.429 ;
        RECT  1.026 38.871 58.104 38.889 ;
        RECT  1.026 38.331 58.104 38.349 ;
        RECT  1.026 37.791 58.104 37.809 ;
        RECT  1.026 37.251 58.104 37.269 ;
        RECT  1.026 36.711 58.104 36.729 ;
        RECT  1.026 36.171 58.104 36.189 ;
        RECT  1.026 35.631 58.104 35.649 ;
        RECT  1.026 35.091 58.104 35.109 ;
        RECT  1.026 34.551 58.104 34.569 ;
        RECT  1.026 34.011 58.104 34.029 ;
        RECT  1.026 33.471 58.104 33.489 ;
        RECT  1.026 32.931 58.104 32.949 ;
        RECT  1.026 32.391 58.104 32.409 ;
        RECT  1.026 31.851 58.104 31.869 ;
        RECT  1.026 31.311 58.104 31.329 ;
        RECT  1.026 30.771 58.104 30.789 ;
        RECT  1.026 30.231 58.104 30.249 ;
        RECT  1.026 29.691 58.104 29.709 ;
        RECT  1.026 29.151 58.104 29.169 ;
        RECT  1.026 28.611 58.104 28.629 ;
        RECT  1.026 28.071 58.104 28.089 ;
        RECT  1.026 27.531 58.104 27.549 ;
        RECT  1.026 26.991 58.104 27.009 ;
        RECT  1.026 26.451 58.104 26.469 ;
        RECT  1.026 25.911 58.104 25.929 ;
        RECT  1.026 25.371 58.104 25.389 ;
        RECT  1.026 24.831 58.104 24.849 ;
        RECT  1.026 24.291 58.104 24.309 ;
        RECT  1.026 23.751 58.104 23.769 ;
        RECT  1.026 23.211 58.104 23.229 ;
        RECT  1.026 22.671 58.104 22.689 ;
        RECT  1.026 22.131 58.104 22.149 ;
        RECT  1.026 21.591 58.104 21.609 ;
        RECT  1.026 21.051 58.104 21.069 ;
        RECT  1.026 20.511 58.104 20.529 ;
        RECT  1.026 19.971 58.104 19.989 ;
        RECT  1.026 19.431 58.104 19.449 ;
        RECT  1.026 18.891 58.104 18.909 ;
        RECT  1.026 18.351 58.104 18.369 ;
        RECT  1.026 17.811 58.104 17.829 ;
        RECT  1.026 17.271 58.104 17.289 ;
        RECT  1.026 16.731 58.104 16.749 ;
        RECT  1.026 16.191 58.104 16.209 ;
        RECT  1.026 15.651 58.104 15.669 ;
        RECT  1.026 15.111 58.104 15.129 ;
        RECT  1.026 14.571 58.104 14.589 ;
        RECT  1.026 14.031 58.104 14.049 ;
        RECT  1.026 13.491 58.104 13.509 ;
        RECT  1.026 12.951 58.104 12.969 ;
        RECT  1.026 12.411 58.104 12.429 ;
        RECT  1.026 11.871 58.104 11.889 ;
        RECT  1.026 11.331 58.104 11.349 ;
        RECT  1.026 10.791 58.104 10.809 ;
        RECT  1.026 10.251 58.104 10.269 ;
        RECT  1.026 9.711 58.104 9.729 ;
        RECT  1.026 9.171 58.104 9.189 ;
        RECT  1.026 8.631 58.104 8.649 ;
        RECT  1.026 8.091 58.104 8.109 ;
        RECT  1.026 7.551 58.104 7.569 ;
        RECT  1.026 7.011 58.104 7.029 ;
        RECT  1.026 6.471 58.104 6.489 ;
        RECT  1.026 5.931 58.104 5.949 ;
        RECT  1.026 5.391 58.104 5.409 ;
        RECT  1.026 4.851 58.104 4.869 ;
        RECT  1.026 4.311 58.104 4.329 ;
        RECT  1.026 3.771 58.104 3.789 ;
        RECT  1.026 3.231 58.104 3.249 ;
        RECT  1.026 2.691 58.104 2.709 ;
        RECT  1.026 2.151 58.104 2.169 ;
        RECT  1.026 1.611 58.104 1.629 ;
        RECT  1.026 1.071 58.104 1.089 ;
      VIA 54.462 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 48.558 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 42.654 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 55.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 49.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 43.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 54.462 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 57.763 54.507 57.797 ;
      VIA 54.462 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 57.223 54.507 57.257 ;
      VIA 54.462 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 56.683 54.507 56.717 ;
      VIA 54.462 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 56.143 54.507 56.177 ;
      VIA 54.462 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 55.603 54.507 55.637 ;
      VIA 54.462 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 55.063 54.507 55.097 ;
      VIA 54.462 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 54.523 54.507 54.557 ;
      VIA 54.462 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 53.983 54.507 54.017 ;
      VIA 54.462 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 53.443 54.507 53.477 ;
      VIA 54.462 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 52.903 54.507 52.937 ;
      VIA 54.462 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 52.363 54.507 52.397 ;
      VIA 54.462 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 51.823 54.507 51.857 ;
      VIA 54.462 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 51.283 54.507 51.317 ;
      VIA 54.462 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 50.743 54.507 50.777 ;
      VIA 54.462 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 50.203 54.507 50.237 ;
      VIA 54.462 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 49.663 54.507 49.697 ;
      VIA 54.462 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 49.123 54.507 49.157 ;
      VIA 54.462 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 48.583 54.507 48.617 ;
      VIA 54.462 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 48.043 54.507 48.077 ;
      VIA 54.462 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 47.503 54.507 47.537 ;
      VIA 54.462 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 46.963 54.507 46.997 ;
      VIA 54.462 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 46.423 54.507 46.457 ;
      VIA 54.462 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 45.883 54.507 45.917 ;
      VIA 54.462 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 45.343 54.507 45.377 ;
      VIA 54.462 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 44.803 54.507 44.837 ;
      VIA 54.462 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 44.263 54.507 44.297 ;
      VIA 54.462 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 43.723 54.507 43.757 ;
      VIA 54.462 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 43.183 54.507 43.217 ;
      VIA 54.462 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 42.643 54.507 42.677 ;
      VIA 54.462 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 42.103 54.507 42.137 ;
      VIA 54.462 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 41.563 54.507 41.597 ;
      VIA 54.462 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 41.023 54.507 41.057 ;
      VIA 54.462 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 40.483 54.507 40.517 ;
      VIA 54.462 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 39.943 54.507 39.977 ;
      VIA 54.462 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 39.403 54.507 39.437 ;
      VIA 54.462 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 38.863 54.507 38.897 ;
      VIA 54.462 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 38.323 54.507 38.357 ;
      VIA 54.462 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 37.783 54.507 37.817 ;
      VIA 54.462 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 37.243 54.507 37.277 ;
      VIA 54.462 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 36.703 54.507 36.737 ;
      VIA 54.462 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 36.163 54.507 36.197 ;
      VIA 54.462 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 35.623 54.507 35.657 ;
      VIA 54.462 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 35.083 54.507 35.117 ;
      VIA 54.462 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 34.543 54.507 34.577 ;
      VIA 54.462 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 34.003 54.507 34.037 ;
      VIA 54.462 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 33.463 54.507 33.497 ;
      VIA 54.462 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 32.923 54.507 32.957 ;
      VIA 54.462 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 32.383 54.507 32.417 ;
      VIA 54.462 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 31.843 54.507 31.877 ;
      VIA 54.462 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 31.303 54.507 31.337 ;
      VIA 54.462 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 30.763 54.507 30.797 ;
      VIA 54.462 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 30.223 54.507 30.257 ;
      VIA 54.462 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 29.683 54.507 29.717 ;
      VIA 54.462 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 29.143 54.507 29.177 ;
      VIA 54.462 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 28.603 54.507 28.637 ;
      VIA 54.462 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 28.063 54.507 28.097 ;
      VIA 54.462 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 27.523 54.507 27.557 ;
      VIA 54.462 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 26.983 54.507 27.017 ;
      VIA 54.462 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 26.443 54.507 26.477 ;
      VIA 54.462 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 25.903 54.507 25.937 ;
      VIA 54.462 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 25.363 54.507 25.397 ;
      VIA 54.462 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 24.823 54.507 24.857 ;
      VIA 54.462 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 24.283 54.507 24.317 ;
      VIA 54.462 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 23.743 54.507 23.777 ;
      VIA 54.462 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 23.203 54.507 23.237 ;
      VIA 54.462 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 22.663 54.507 22.697 ;
      VIA 54.462 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 22.123 54.507 22.157 ;
      VIA 54.462 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 21.583 54.507 21.617 ;
      VIA 54.462 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 21.043 54.507 21.077 ;
      VIA 54.462 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 20.503 54.507 20.537 ;
      VIA 54.462 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 19.963 54.507 19.997 ;
      VIA 54.462 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 19.423 54.507 19.457 ;
      VIA 54.462 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 18.883 54.507 18.917 ;
      VIA 54.462 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 18.343 54.507 18.377 ;
      VIA 54.462 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 17.803 54.507 17.837 ;
      VIA 54.462 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 17.263 54.507 17.297 ;
      VIA 54.462 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 16.723 54.507 16.757 ;
      VIA 54.462 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 16.183 54.507 16.217 ;
      VIA 54.462 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 15.643 54.507 15.677 ;
      VIA 54.462 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 15.103 54.507 15.137 ;
      VIA 54.462 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 14.563 54.507 14.597 ;
      VIA 54.462 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 14.023 54.507 14.057 ;
      VIA 54.462 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 13.483 54.507 13.517 ;
      VIA 54.462 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 12.943 54.507 12.977 ;
      VIA 54.462 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 12.403 54.507 12.437 ;
      VIA 54.462 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 11.863 54.507 11.897 ;
      VIA 54.462 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 11.323 54.507 11.357 ;
      VIA 54.462 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 10.783 54.507 10.817 ;
      VIA 54.462 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 10.243 54.507 10.277 ;
      VIA 54.462 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 9.703 54.507 9.737 ;
      VIA 54.462 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 9.163 54.507 9.197 ;
      VIA 54.462 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 8.623 54.507 8.657 ;
      VIA 54.462 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 8.083 54.507 8.117 ;
      VIA 54.462 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 7.543 54.507 7.577 ;
      VIA 54.462 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 7.003 54.507 7.037 ;
      VIA 54.462 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 6.463 54.507 6.497 ;
      VIA 54.462 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 5.923 54.507 5.957 ;
      VIA 54.462 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 5.383 54.507 5.417 ;
      VIA 54.462 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 4.843 54.507 4.877 ;
      VIA 54.462 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 4.303 54.507 4.337 ;
      VIA 54.462 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 3.763 54.507 3.797 ;
      VIA 54.462 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 3.223 54.507 3.257 ;
      VIA 54.462 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 2.683 54.507 2.717 ;
      VIA 54.462 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 2.143 54.507 2.177 ;
      VIA 54.462 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 1.603 54.507 1.637 ;
      VIA 54.462 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 54.462 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  54.417 1.063 54.507 1.097 ;
      VIA 54.462 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 54.462 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 57.763 48.603 57.797 ;
      VIA 48.558 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 57.223 48.603 57.257 ;
      VIA 48.558 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 56.683 48.603 56.717 ;
      VIA 48.558 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 56.143 48.603 56.177 ;
      VIA 48.558 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 55.603 48.603 55.637 ;
      VIA 48.558 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 55.063 48.603 55.097 ;
      VIA 48.558 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 54.523 48.603 54.557 ;
      VIA 48.558 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 53.983 48.603 54.017 ;
      VIA 48.558 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 53.443 48.603 53.477 ;
      VIA 48.558 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 52.903 48.603 52.937 ;
      VIA 48.558 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 52.363 48.603 52.397 ;
      VIA 48.558 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 51.823 48.603 51.857 ;
      VIA 48.558 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 51.283 48.603 51.317 ;
      VIA 48.558 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 50.743 48.603 50.777 ;
      VIA 48.558 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 50.203 48.603 50.237 ;
      VIA 48.558 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 49.663 48.603 49.697 ;
      VIA 48.558 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 49.123 48.603 49.157 ;
      VIA 48.558 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 48.583 48.603 48.617 ;
      VIA 48.558 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 48.043 48.603 48.077 ;
      VIA 48.558 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 47.503 48.603 47.537 ;
      VIA 48.558 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 46.963 48.603 46.997 ;
      VIA 48.558 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 46.423 48.603 46.457 ;
      VIA 48.558 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 45.883 48.603 45.917 ;
      VIA 48.558 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 45.343 48.603 45.377 ;
      VIA 48.558 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 44.803 48.603 44.837 ;
      VIA 48.558 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 44.263 48.603 44.297 ;
      VIA 48.558 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 43.723 48.603 43.757 ;
      VIA 48.558 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 43.183 48.603 43.217 ;
      VIA 48.558 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 42.643 48.603 42.677 ;
      VIA 48.558 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 42.103 48.603 42.137 ;
      VIA 48.558 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 41.563 48.603 41.597 ;
      VIA 48.558 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 41.023 48.603 41.057 ;
      VIA 48.558 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 40.483 48.603 40.517 ;
      VIA 48.558 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 39.943 48.603 39.977 ;
      VIA 48.558 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 39.403 48.603 39.437 ;
      VIA 48.558 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 38.863 48.603 38.897 ;
      VIA 48.558 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 38.323 48.603 38.357 ;
      VIA 48.558 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 37.783 48.603 37.817 ;
      VIA 48.558 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 37.243 48.603 37.277 ;
      VIA 48.558 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 36.703 48.603 36.737 ;
      VIA 48.558 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 36.163 48.603 36.197 ;
      VIA 48.558 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 35.623 48.603 35.657 ;
      VIA 48.558 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 35.083 48.603 35.117 ;
      VIA 48.558 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 34.543 48.603 34.577 ;
      VIA 48.558 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 34.003 48.603 34.037 ;
      VIA 48.558 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 33.463 48.603 33.497 ;
      VIA 48.558 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 32.923 48.603 32.957 ;
      VIA 48.558 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 32.383 48.603 32.417 ;
      VIA 48.558 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 31.843 48.603 31.877 ;
      VIA 48.558 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 31.303 48.603 31.337 ;
      VIA 48.558 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 30.763 48.603 30.797 ;
      VIA 48.558 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 30.223 48.603 30.257 ;
      VIA 48.558 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 29.683 48.603 29.717 ;
      VIA 48.558 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 29.143 48.603 29.177 ;
      VIA 48.558 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 28.603 48.603 28.637 ;
      VIA 48.558 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 28.063 48.603 28.097 ;
      VIA 48.558 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 27.523 48.603 27.557 ;
      VIA 48.558 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 26.983 48.603 27.017 ;
      VIA 48.558 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 26.443 48.603 26.477 ;
      VIA 48.558 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 25.903 48.603 25.937 ;
      VIA 48.558 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 25.363 48.603 25.397 ;
      VIA 48.558 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 24.823 48.603 24.857 ;
      VIA 48.558 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 24.283 48.603 24.317 ;
      VIA 48.558 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 23.743 48.603 23.777 ;
      VIA 48.558 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 23.203 48.603 23.237 ;
      VIA 48.558 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 22.663 48.603 22.697 ;
      VIA 48.558 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 22.123 48.603 22.157 ;
      VIA 48.558 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 21.583 48.603 21.617 ;
      VIA 48.558 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 21.043 48.603 21.077 ;
      VIA 48.558 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 20.503 48.603 20.537 ;
      VIA 48.558 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 19.963 48.603 19.997 ;
      VIA 48.558 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 19.423 48.603 19.457 ;
      VIA 48.558 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 18.883 48.603 18.917 ;
      VIA 48.558 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 18.343 48.603 18.377 ;
      VIA 48.558 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 17.803 48.603 17.837 ;
      VIA 48.558 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 17.263 48.603 17.297 ;
      VIA 48.558 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 16.723 48.603 16.757 ;
      VIA 48.558 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 16.183 48.603 16.217 ;
      VIA 48.558 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 15.643 48.603 15.677 ;
      VIA 48.558 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 15.103 48.603 15.137 ;
      VIA 48.558 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 14.563 48.603 14.597 ;
      VIA 48.558 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 14.023 48.603 14.057 ;
      VIA 48.558 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 13.483 48.603 13.517 ;
      VIA 48.558 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 12.943 48.603 12.977 ;
      VIA 48.558 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 12.403 48.603 12.437 ;
      VIA 48.558 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 11.863 48.603 11.897 ;
      VIA 48.558 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 11.323 48.603 11.357 ;
      VIA 48.558 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 10.783 48.603 10.817 ;
      VIA 48.558 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 10.243 48.603 10.277 ;
      VIA 48.558 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 9.703 48.603 9.737 ;
      VIA 48.558 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 9.163 48.603 9.197 ;
      VIA 48.558 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 8.623 48.603 8.657 ;
      VIA 48.558 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 8.083 48.603 8.117 ;
      VIA 48.558 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 7.543 48.603 7.577 ;
      VIA 48.558 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 7.003 48.603 7.037 ;
      VIA 48.558 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 6.463 48.603 6.497 ;
      VIA 48.558 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 5.923 48.603 5.957 ;
      VIA 48.558 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 5.383 48.603 5.417 ;
      VIA 48.558 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 4.843 48.603 4.877 ;
      VIA 48.558 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 4.303 48.603 4.337 ;
      VIA 48.558 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 3.763 48.603 3.797 ;
      VIA 48.558 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 3.223 48.603 3.257 ;
      VIA 48.558 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 2.683 48.603 2.717 ;
      VIA 48.558 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 2.143 48.603 2.177 ;
      VIA 48.558 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 1.603 48.603 1.637 ;
      VIA 48.558 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 48.558 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  48.513 1.063 48.603 1.097 ;
      VIA 48.558 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 48.558 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 57.763 42.699 57.797 ;
      VIA 42.654 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 57.223 42.699 57.257 ;
      VIA 42.654 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 56.683 42.699 56.717 ;
      VIA 42.654 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 56.143 42.699 56.177 ;
      VIA 42.654 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 55.603 42.699 55.637 ;
      VIA 42.654 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 55.063 42.699 55.097 ;
      VIA 42.654 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 54.523 42.699 54.557 ;
      VIA 42.654 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 53.983 42.699 54.017 ;
      VIA 42.654 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 53.443 42.699 53.477 ;
      VIA 42.654 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 52.903 42.699 52.937 ;
      VIA 42.654 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 52.363 42.699 52.397 ;
      VIA 42.654 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 51.823 42.699 51.857 ;
      VIA 42.654 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 51.283 42.699 51.317 ;
      VIA 42.654 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 50.743 42.699 50.777 ;
      VIA 42.654 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 50.203 42.699 50.237 ;
      VIA 42.654 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 49.663 42.699 49.697 ;
      VIA 42.654 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 49.123 42.699 49.157 ;
      VIA 42.654 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 48.583 42.699 48.617 ;
      VIA 42.654 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 48.043 42.699 48.077 ;
      VIA 42.654 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 47.503 42.699 47.537 ;
      VIA 42.654 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 46.963 42.699 46.997 ;
      VIA 42.654 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 46.423 42.699 46.457 ;
      VIA 42.654 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 45.883 42.699 45.917 ;
      VIA 42.654 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 45.343 42.699 45.377 ;
      VIA 42.654 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 44.803 42.699 44.837 ;
      VIA 42.654 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 44.263 42.699 44.297 ;
      VIA 42.654 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 43.723 42.699 43.757 ;
      VIA 42.654 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 43.183 42.699 43.217 ;
      VIA 42.654 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 42.643 42.699 42.677 ;
      VIA 42.654 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 42.103 42.699 42.137 ;
      VIA 42.654 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 41.563 42.699 41.597 ;
      VIA 42.654 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 41.023 42.699 41.057 ;
      VIA 42.654 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 40.483 42.699 40.517 ;
      VIA 42.654 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 39.943 42.699 39.977 ;
      VIA 42.654 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 39.403 42.699 39.437 ;
      VIA 42.654 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 38.863 42.699 38.897 ;
      VIA 42.654 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 38.323 42.699 38.357 ;
      VIA 42.654 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 37.783 42.699 37.817 ;
      VIA 42.654 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 37.243 42.699 37.277 ;
      VIA 42.654 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 36.703 42.699 36.737 ;
      VIA 42.654 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 36.163 42.699 36.197 ;
      VIA 42.654 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 35.623 42.699 35.657 ;
      VIA 42.654 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 35.083 42.699 35.117 ;
      VIA 42.654 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 34.543 42.699 34.577 ;
      VIA 42.654 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 34.003 42.699 34.037 ;
      VIA 42.654 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 33.463 42.699 33.497 ;
      VIA 42.654 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 32.923 42.699 32.957 ;
      VIA 42.654 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 32.383 42.699 32.417 ;
      VIA 42.654 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 31.843 42.699 31.877 ;
      VIA 42.654 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 31.303 42.699 31.337 ;
      VIA 42.654 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 30.763 42.699 30.797 ;
      VIA 42.654 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 30.223 42.699 30.257 ;
      VIA 42.654 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 29.683 42.699 29.717 ;
      VIA 42.654 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 29.143 42.699 29.177 ;
      VIA 42.654 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 28.603 42.699 28.637 ;
      VIA 42.654 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 28.063 42.699 28.097 ;
      VIA 42.654 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 27.523 42.699 27.557 ;
      VIA 42.654 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 26.983 42.699 27.017 ;
      VIA 42.654 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 26.443 42.699 26.477 ;
      VIA 42.654 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 25.903 42.699 25.937 ;
      VIA 42.654 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 25.363 42.699 25.397 ;
      VIA 42.654 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 24.823 42.699 24.857 ;
      VIA 42.654 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 24.283 42.699 24.317 ;
      VIA 42.654 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 23.743 42.699 23.777 ;
      VIA 42.654 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 23.203 42.699 23.237 ;
      VIA 42.654 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 22.663 42.699 22.697 ;
      VIA 42.654 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 22.123 42.699 22.157 ;
      VIA 42.654 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 21.583 42.699 21.617 ;
      VIA 42.654 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 21.043 42.699 21.077 ;
      VIA 42.654 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 20.503 42.699 20.537 ;
      VIA 42.654 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 19.963 42.699 19.997 ;
      VIA 42.654 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 19.423 42.699 19.457 ;
      VIA 42.654 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 18.883 42.699 18.917 ;
      VIA 42.654 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 18.343 42.699 18.377 ;
      VIA 42.654 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 17.803 42.699 17.837 ;
      VIA 42.654 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 17.263 42.699 17.297 ;
      VIA 42.654 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 16.723 42.699 16.757 ;
      VIA 42.654 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 16.183 42.699 16.217 ;
      VIA 42.654 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 15.643 42.699 15.677 ;
      VIA 42.654 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 15.103 42.699 15.137 ;
      VIA 42.654 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 14.563 42.699 14.597 ;
      VIA 42.654 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 14.023 42.699 14.057 ;
      VIA 42.654 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 13.483 42.699 13.517 ;
      VIA 42.654 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 12.943 42.699 12.977 ;
      VIA 42.654 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 12.403 42.699 12.437 ;
      VIA 42.654 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 11.863 42.699 11.897 ;
      VIA 42.654 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 11.323 42.699 11.357 ;
      VIA 42.654 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 10.783 42.699 10.817 ;
      VIA 42.654 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 10.243 42.699 10.277 ;
      VIA 42.654 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 9.703 42.699 9.737 ;
      VIA 42.654 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 9.163 42.699 9.197 ;
      VIA 42.654 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 8.623 42.699 8.657 ;
      VIA 42.654 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 8.083 42.699 8.117 ;
      VIA 42.654 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 7.543 42.699 7.577 ;
      VIA 42.654 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 7.003 42.699 7.037 ;
      VIA 42.654 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 6.463 42.699 6.497 ;
      VIA 42.654 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 5.923 42.699 5.957 ;
      VIA 42.654 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 5.383 42.699 5.417 ;
      VIA 42.654 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 4.843 42.699 4.877 ;
      VIA 42.654 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 4.303 42.699 4.337 ;
      VIA 42.654 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 3.763 42.699 3.797 ;
      VIA 42.654 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 3.223 42.699 3.257 ;
      VIA 42.654 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 2.683 42.699 2.717 ;
      VIA 42.654 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 2.143 42.699 2.177 ;
      VIA 42.654 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 1.603 42.699 1.637 ;
      VIA 42.654 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 42.654 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  42.609 1.063 42.699 1.097 ;
      VIA 42.654 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 42.654 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 57.763 36.795 57.797 ;
      VIA 36.75 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 57.223 36.795 57.257 ;
      VIA 36.75 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 56.683 36.795 56.717 ;
      VIA 36.75 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 56.143 36.795 56.177 ;
      VIA 36.75 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 55.603 36.795 55.637 ;
      VIA 36.75 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 55.063 36.795 55.097 ;
      VIA 36.75 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 54.523 36.795 54.557 ;
      VIA 36.75 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 53.983 36.795 54.017 ;
      VIA 36.75 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 53.443 36.795 53.477 ;
      VIA 36.75 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 52.903 36.795 52.937 ;
      VIA 36.75 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 52.363 36.795 52.397 ;
      VIA 36.75 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 51.823 36.795 51.857 ;
      VIA 36.75 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 51.283 36.795 51.317 ;
      VIA 36.75 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 50.743 36.795 50.777 ;
      VIA 36.75 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 50.203 36.795 50.237 ;
      VIA 36.75 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 49.663 36.795 49.697 ;
      VIA 36.75 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 49.123 36.795 49.157 ;
      VIA 36.75 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 48.583 36.795 48.617 ;
      VIA 36.75 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 48.043 36.795 48.077 ;
      VIA 36.75 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 47.503 36.795 47.537 ;
      VIA 36.75 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 46.963 36.795 46.997 ;
      VIA 36.75 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 46.423 36.795 46.457 ;
      VIA 36.75 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 45.883 36.795 45.917 ;
      VIA 36.75 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 45.343 36.795 45.377 ;
      VIA 36.75 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 44.803 36.795 44.837 ;
      VIA 36.75 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 44.263 36.795 44.297 ;
      VIA 36.75 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 43.723 36.795 43.757 ;
      VIA 36.75 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 43.183 36.795 43.217 ;
      VIA 36.75 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 42.643 36.795 42.677 ;
      VIA 36.75 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 42.103 36.795 42.137 ;
      VIA 36.75 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 41.563 36.795 41.597 ;
      VIA 36.75 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 41.023 36.795 41.057 ;
      VIA 36.75 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 40.483 36.795 40.517 ;
      VIA 36.75 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.943 36.795 39.977 ;
      VIA 36.75 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.403 36.795 39.437 ;
      VIA 36.75 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.863 36.795 38.897 ;
      VIA 36.75 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.323 36.795 38.357 ;
      VIA 36.75 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.783 36.795 37.817 ;
      VIA 36.75 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.243 36.795 37.277 ;
      VIA 36.75 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.703 36.795 36.737 ;
      VIA 36.75 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.163 36.795 36.197 ;
      VIA 36.75 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.623 36.795 35.657 ;
      VIA 36.75 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.083 36.795 35.117 ;
      VIA 36.75 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.543 36.795 34.577 ;
      VIA 36.75 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.003 36.795 34.037 ;
      VIA 36.75 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 33.463 36.795 33.497 ;
      VIA 36.75 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.923 36.795 32.957 ;
      VIA 36.75 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.383 36.795 32.417 ;
      VIA 36.75 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.843 36.795 31.877 ;
      VIA 36.75 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.303 36.795 31.337 ;
      VIA 36.75 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.763 36.795 30.797 ;
      VIA 36.75 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.223 36.795 30.257 ;
      VIA 36.75 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.683 36.795 29.717 ;
      VIA 36.75 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.143 36.795 29.177 ;
      VIA 36.75 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.603 36.795 28.637 ;
      VIA 36.75 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.063 36.795 28.097 ;
      VIA 36.75 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 27.523 36.795 27.557 ;
      VIA 36.75 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.983 36.795 27.017 ;
      VIA 36.75 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.443 36.795 26.477 ;
      VIA 36.75 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.903 36.795 25.937 ;
      VIA 36.75 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.363 36.795 25.397 ;
      VIA 36.75 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.823 36.795 24.857 ;
      VIA 36.75 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.283 36.795 24.317 ;
      VIA 36.75 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.743 36.795 23.777 ;
      VIA 36.75 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.203 36.795 23.237 ;
      VIA 36.75 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.663 36.795 22.697 ;
      VIA 36.75 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.123 36.795 22.157 ;
      VIA 36.75 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.583 36.795 21.617 ;
      VIA 36.75 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.043 36.795 21.077 ;
      VIA 36.75 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 20.503 36.795 20.537 ;
      VIA 36.75 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.963 36.795 19.997 ;
      VIA 36.75 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.423 36.795 19.457 ;
      VIA 36.75 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.883 36.795 18.917 ;
      VIA 36.75 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.343 36.795 18.377 ;
      VIA 36.75 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.803 36.795 17.837 ;
      VIA 36.75 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.263 36.795 17.297 ;
      VIA 36.75 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.723 36.795 16.757 ;
      VIA 36.75 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.183 36.795 16.217 ;
      VIA 36.75 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.643 36.795 15.677 ;
      VIA 36.75 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.103 36.795 15.137 ;
      VIA 36.75 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.563 36.795 14.597 ;
      VIA 36.75 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.023 36.795 14.057 ;
      VIA 36.75 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 13.483 36.795 13.517 ;
      VIA 36.75 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.943 36.795 12.977 ;
      VIA 36.75 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.403 36.795 12.437 ;
      VIA 36.75 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.863 36.795 11.897 ;
      VIA 36.75 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.323 36.795 11.357 ;
      VIA 36.75 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.783 36.795 10.817 ;
      VIA 36.75 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.243 36.795 10.277 ;
      VIA 36.75 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.703 36.795 9.737 ;
      VIA 36.75 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.163 36.795 9.197 ;
      VIA 36.75 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.623 36.795 8.657 ;
      VIA 36.75 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.083 36.795 8.117 ;
      VIA 36.75 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.543 36.795 7.577 ;
      VIA 36.75 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.003 36.795 7.037 ;
      VIA 36.75 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 6.463 36.795 6.497 ;
      VIA 36.75 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.923 36.795 5.957 ;
      VIA 36.75 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.383 36.795 5.417 ;
      VIA 36.75 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.843 36.795 4.877 ;
      VIA 36.75 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.303 36.795 4.337 ;
      VIA 36.75 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.763 36.795 3.797 ;
      VIA 36.75 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.223 36.795 3.257 ;
      VIA 36.75 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.683 36.795 2.717 ;
      VIA 36.75 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.143 36.795 2.177 ;
      VIA 36.75 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.603 36.795 1.637 ;
      VIA 36.75 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.063 36.795 1.097 ;
      VIA 36.75 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 57.763 30.891 57.797 ;
      VIA 30.846 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 57.223 30.891 57.257 ;
      VIA 30.846 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 56.683 30.891 56.717 ;
      VIA 30.846 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 56.143 30.891 56.177 ;
      VIA 30.846 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 55.603 30.891 55.637 ;
      VIA 30.846 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 55.063 30.891 55.097 ;
      VIA 30.846 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 54.523 30.891 54.557 ;
      VIA 30.846 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 53.983 30.891 54.017 ;
      VIA 30.846 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 53.443 30.891 53.477 ;
      VIA 30.846 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 52.903 30.891 52.937 ;
      VIA 30.846 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 52.363 30.891 52.397 ;
      VIA 30.846 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 51.823 30.891 51.857 ;
      VIA 30.846 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 51.283 30.891 51.317 ;
      VIA 30.846 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 50.743 30.891 50.777 ;
      VIA 30.846 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 50.203 30.891 50.237 ;
      VIA 30.846 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 49.663 30.891 49.697 ;
      VIA 30.846 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 49.123 30.891 49.157 ;
      VIA 30.846 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 48.583 30.891 48.617 ;
      VIA 30.846 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 48.043 30.891 48.077 ;
      VIA 30.846 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 47.503 30.891 47.537 ;
      VIA 30.846 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 46.963 30.891 46.997 ;
      VIA 30.846 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 46.423 30.891 46.457 ;
      VIA 30.846 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 45.883 30.891 45.917 ;
      VIA 30.846 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 45.343 30.891 45.377 ;
      VIA 30.846 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 44.803 30.891 44.837 ;
      VIA 30.846 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 44.263 30.891 44.297 ;
      VIA 30.846 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 43.723 30.891 43.757 ;
      VIA 30.846 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 43.183 30.891 43.217 ;
      VIA 30.846 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 42.643 30.891 42.677 ;
      VIA 30.846 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 42.103 30.891 42.137 ;
      VIA 30.846 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 41.563 30.891 41.597 ;
      VIA 30.846 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 41.023 30.891 41.057 ;
      VIA 30.846 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 40.483 30.891 40.517 ;
      VIA 30.846 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.943 30.891 39.977 ;
      VIA 30.846 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.403 30.891 39.437 ;
      VIA 30.846 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.863 30.891 38.897 ;
      VIA 30.846 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.323 30.891 38.357 ;
      VIA 30.846 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.783 30.891 37.817 ;
      VIA 30.846 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.243 30.891 37.277 ;
      VIA 30.846 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.703 30.891 36.737 ;
      VIA 30.846 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.163 30.891 36.197 ;
      VIA 30.846 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.623 30.891 35.657 ;
      VIA 30.846 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.083 30.891 35.117 ;
      VIA 30.846 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.543 30.891 34.577 ;
      VIA 30.846 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.003 30.891 34.037 ;
      VIA 30.846 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 33.463 30.891 33.497 ;
      VIA 30.846 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.923 30.891 32.957 ;
      VIA 30.846 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.383 30.891 32.417 ;
      VIA 30.846 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.843 30.891 31.877 ;
      VIA 30.846 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.303 30.891 31.337 ;
      VIA 30.846 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.763 30.891 30.797 ;
      VIA 30.846 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.223 30.891 30.257 ;
      VIA 30.846 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.683 30.891 29.717 ;
      VIA 30.846 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.143 30.891 29.177 ;
      VIA 30.846 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.603 30.891 28.637 ;
      VIA 30.846 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.063 30.891 28.097 ;
      VIA 30.846 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 27.523 30.891 27.557 ;
      VIA 30.846 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.983 30.891 27.017 ;
      VIA 30.846 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.443 30.891 26.477 ;
      VIA 30.846 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.903 30.891 25.937 ;
      VIA 30.846 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.363 30.891 25.397 ;
      VIA 30.846 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.823 30.891 24.857 ;
      VIA 30.846 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.283 30.891 24.317 ;
      VIA 30.846 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.743 30.891 23.777 ;
      VIA 30.846 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.203 30.891 23.237 ;
      VIA 30.846 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.663 30.891 22.697 ;
      VIA 30.846 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.123 30.891 22.157 ;
      VIA 30.846 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.583 30.891 21.617 ;
      VIA 30.846 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.043 30.891 21.077 ;
      VIA 30.846 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 20.503 30.891 20.537 ;
      VIA 30.846 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.963 30.891 19.997 ;
      VIA 30.846 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.423 30.891 19.457 ;
      VIA 30.846 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.883 30.891 18.917 ;
      VIA 30.846 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.343 30.891 18.377 ;
      VIA 30.846 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.803 30.891 17.837 ;
      VIA 30.846 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.263 30.891 17.297 ;
      VIA 30.846 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.723 30.891 16.757 ;
      VIA 30.846 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.183 30.891 16.217 ;
      VIA 30.846 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.643 30.891 15.677 ;
      VIA 30.846 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.103 30.891 15.137 ;
      VIA 30.846 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.563 30.891 14.597 ;
      VIA 30.846 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.023 30.891 14.057 ;
      VIA 30.846 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 13.483 30.891 13.517 ;
      VIA 30.846 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.943 30.891 12.977 ;
      VIA 30.846 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.403 30.891 12.437 ;
      VIA 30.846 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.863 30.891 11.897 ;
      VIA 30.846 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.323 30.891 11.357 ;
      VIA 30.846 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.783 30.891 10.817 ;
      VIA 30.846 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.243 30.891 10.277 ;
      VIA 30.846 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.703 30.891 9.737 ;
      VIA 30.846 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.163 30.891 9.197 ;
      VIA 30.846 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.623 30.891 8.657 ;
      VIA 30.846 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.083 30.891 8.117 ;
      VIA 30.846 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.543 30.891 7.577 ;
      VIA 30.846 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.003 30.891 7.037 ;
      VIA 30.846 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 6.463 30.891 6.497 ;
      VIA 30.846 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.923 30.891 5.957 ;
      VIA 30.846 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.383 30.891 5.417 ;
      VIA 30.846 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.843 30.891 4.877 ;
      VIA 30.846 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.303 30.891 4.337 ;
      VIA 30.846 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.763 30.891 3.797 ;
      VIA 30.846 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.223 30.891 3.257 ;
      VIA 30.846 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.683 30.891 2.717 ;
      VIA 30.846 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.143 30.891 2.177 ;
      VIA 30.846 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.603 30.891 1.637 ;
      VIA 30.846 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.063 30.891 1.097 ;
      VIA 30.846 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 57.763 24.987 57.797 ;
      VIA 24.942 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 57.223 24.987 57.257 ;
      VIA 24.942 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 56.683 24.987 56.717 ;
      VIA 24.942 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 56.143 24.987 56.177 ;
      VIA 24.942 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 55.603 24.987 55.637 ;
      VIA 24.942 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 55.063 24.987 55.097 ;
      VIA 24.942 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 54.523 24.987 54.557 ;
      VIA 24.942 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 53.983 24.987 54.017 ;
      VIA 24.942 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 53.443 24.987 53.477 ;
      VIA 24.942 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 52.903 24.987 52.937 ;
      VIA 24.942 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 52.363 24.987 52.397 ;
      VIA 24.942 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 51.823 24.987 51.857 ;
      VIA 24.942 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 51.283 24.987 51.317 ;
      VIA 24.942 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 50.743 24.987 50.777 ;
      VIA 24.942 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 50.203 24.987 50.237 ;
      VIA 24.942 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 49.663 24.987 49.697 ;
      VIA 24.942 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 49.123 24.987 49.157 ;
      VIA 24.942 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 48.583 24.987 48.617 ;
      VIA 24.942 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 48.043 24.987 48.077 ;
      VIA 24.942 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 47.503 24.987 47.537 ;
      VIA 24.942 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 46.963 24.987 46.997 ;
      VIA 24.942 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 46.423 24.987 46.457 ;
      VIA 24.942 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 45.883 24.987 45.917 ;
      VIA 24.942 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 45.343 24.987 45.377 ;
      VIA 24.942 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 44.803 24.987 44.837 ;
      VIA 24.942 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 44.263 24.987 44.297 ;
      VIA 24.942 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 43.723 24.987 43.757 ;
      VIA 24.942 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 43.183 24.987 43.217 ;
      VIA 24.942 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 42.643 24.987 42.677 ;
      VIA 24.942 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 42.103 24.987 42.137 ;
      VIA 24.942 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 41.563 24.987 41.597 ;
      VIA 24.942 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 41.023 24.987 41.057 ;
      VIA 24.942 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 40.483 24.987 40.517 ;
      VIA 24.942 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.943 24.987 39.977 ;
      VIA 24.942 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.403 24.987 39.437 ;
      VIA 24.942 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.863 24.987 38.897 ;
      VIA 24.942 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.323 24.987 38.357 ;
      VIA 24.942 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.783 24.987 37.817 ;
      VIA 24.942 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.243 24.987 37.277 ;
      VIA 24.942 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.703 24.987 36.737 ;
      VIA 24.942 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.163 24.987 36.197 ;
      VIA 24.942 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.623 24.987 35.657 ;
      VIA 24.942 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.083 24.987 35.117 ;
      VIA 24.942 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.543 24.987 34.577 ;
      VIA 24.942 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.003 24.987 34.037 ;
      VIA 24.942 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 33.463 24.987 33.497 ;
      VIA 24.942 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.923 24.987 32.957 ;
      VIA 24.942 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.383 24.987 32.417 ;
      VIA 24.942 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.843 24.987 31.877 ;
      VIA 24.942 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.303 24.987 31.337 ;
      VIA 24.942 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.763 24.987 30.797 ;
      VIA 24.942 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.223 24.987 30.257 ;
      VIA 24.942 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.683 24.987 29.717 ;
      VIA 24.942 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.143 24.987 29.177 ;
      VIA 24.942 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.603 24.987 28.637 ;
      VIA 24.942 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.063 24.987 28.097 ;
      VIA 24.942 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 27.523 24.987 27.557 ;
      VIA 24.942 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.983 24.987 27.017 ;
      VIA 24.942 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.443 24.987 26.477 ;
      VIA 24.942 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.903 24.987 25.937 ;
      VIA 24.942 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.363 24.987 25.397 ;
      VIA 24.942 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.823 24.987 24.857 ;
      VIA 24.942 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.283 24.987 24.317 ;
      VIA 24.942 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.743 24.987 23.777 ;
      VIA 24.942 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.203 24.987 23.237 ;
      VIA 24.942 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.663 24.987 22.697 ;
      VIA 24.942 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.123 24.987 22.157 ;
      VIA 24.942 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.583 24.987 21.617 ;
      VIA 24.942 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.043 24.987 21.077 ;
      VIA 24.942 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 20.503 24.987 20.537 ;
      VIA 24.942 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.963 24.987 19.997 ;
      VIA 24.942 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.423 24.987 19.457 ;
      VIA 24.942 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.883 24.987 18.917 ;
      VIA 24.942 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.343 24.987 18.377 ;
      VIA 24.942 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.803 24.987 17.837 ;
      VIA 24.942 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.263 24.987 17.297 ;
      VIA 24.942 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.723 24.987 16.757 ;
      VIA 24.942 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.183 24.987 16.217 ;
      VIA 24.942 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.643 24.987 15.677 ;
      VIA 24.942 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.103 24.987 15.137 ;
      VIA 24.942 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.563 24.987 14.597 ;
      VIA 24.942 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.023 24.987 14.057 ;
      VIA 24.942 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 13.483 24.987 13.517 ;
      VIA 24.942 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.943 24.987 12.977 ;
      VIA 24.942 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.403 24.987 12.437 ;
      VIA 24.942 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.863 24.987 11.897 ;
      VIA 24.942 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.323 24.987 11.357 ;
      VIA 24.942 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.783 24.987 10.817 ;
      VIA 24.942 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.243 24.987 10.277 ;
      VIA 24.942 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.703 24.987 9.737 ;
      VIA 24.942 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.163 24.987 9.197 ;
      VIA 24.942 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.623 24.987 8.657 ;
      VIA 24.942 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.083 24.987 8.117 ;
      VIA 24.942 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.543 24.987 7.577 ;
      VIA 24.942 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.003 24.987 7.037 ;
      VIA 24.942 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 6.463 24.987 6.497 ;
      VIA 24.942 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.923 24.987 5.957 ;
      VIA 24.942 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.383 24.987 5.417 ;
      VIA 24.942 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.843 24.987 4.877 ;
      VIA 24.942 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.303 24.987 4.337 ;
      VIA 24.942 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.763 24.987 3.797 ;
      VIA 24.942 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.223 24.987 3.257 ;
      VIA 24.942 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.683 24.987 2.717 ;
      VIA 24.942 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.143 24.987 2.177 ;
      VIA 24.942 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.603 24.987 1.637 ;
      VIA 24.942 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.063 24.987 1.097 ;
      VIA 24.942 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 57.763 19.083 57.797 ;
      VIA 19.038 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 57.223 19.083 57.257 ;
      VIA 19.038 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 56.683 19.083 56.717 ;
      VIA 19.038 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 56.143 19.083 56.177 ;
      VIA 19.038 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 55.603 19.083 55.637 ;
      VIA 19.038 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 55.063 19.083 55.097 ;
      VIA 19.038 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 54.523 19.083 54.557 ;
      VIA 19.038 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 53.983 19.083 54.017 ;
      VIA 19.038 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 53.443 19.083 53.477 ;
      VIA 19.038 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 52.903 19.083 52.937 ;
      VIA 19.038 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 52.363 19.083 52.397 ;
      VIA 19.038 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 51.823 19.083 51.857 ;
      VIA 19.038 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 51.283 19.083 51.317 ;
      VIA 19.038 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 50.743 19.083 50.777 ;
      VIA 19.038 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 50.203 19.083 50.237 ;
      VIA 19.038 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 49.663 19.083 49.697 ;
      VIA 19.038 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 49.123 19.083 49.157 ;
      VIA 19.038 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 48.583 19.083 48.617 ;
      VIA 19.038 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 48.043 19.083 48.077 ;
      VIA 19.038 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 47.503 19.083 47.537 ;
      VIA 19.038 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 46.963 19.083 46.997 ;
      VIA 19.038 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 46.423 19.083 46.457 ;
      VIA 19.038 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 45.883 19.083 45.917 ;
      VIA 19.038 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 45.343 19.083 45.377 ;
      VIA 19.038 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 44.803 19.083 44.837 ;
      VIA 19.038 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 44.263 19.083 44.297 ;
      VIA 19.038 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 43.723 19.083 43.757 ;
      VIA 19.038 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 43.183 19.083 43.217 ;
      VIA 19.038 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 42.643 19.083 42.677 ;
      VIA 19.038 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 42.103 19.083 42.137 ;
      VIA 19.038 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 41.563 19.083 41.597 ;
      VIA 19.038 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 41.023 19.083 41.057 ;
      VIA 19.038 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 40.483 19.083 40.517 ;
      VIA 19.038 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.943 19.083 39.977 ;
      VIA 19.038 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.403 19.083 39.437 ;
      VIA 19.038 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.863 19.083 38.897 ;
      VIA 19.038 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.323 19.083 38.357 ;
      VIA 19.038 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.783 19.083 37.817 ;
      VIA 19.038 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.243 19.083 37.277 ;
      VIA 19.038 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.703 19.083 36.737 ;
      VIA 19.038 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.163 19.083 36.197 ;
      VIA 19.038 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.623 19.083 35.657 ;
      VIA 19.038 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.083 19.083 35.117 ;
      VIA 19.038 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.543 19.083 34.577 ;
      VIA 19.038 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.003 19.083 34.037 ;
      VIA 19.038 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 33.463 19.083 33.497 ;
      VIA 19.038 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.923 19.083 32.957 ;
      VIA 19.038 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.383 19.083 32.417 ;
      VIA 19.038 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.843 19.083 31.877 ;
      VIA 19.038 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.303 19.083 31.337 ;
      VIA 19.038 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.763 19.083 30.797 ;
      VIA 19.038 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.223 19.083 30.257 ;
      VIA 19.038 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.683 19.083 29.717 ;
      VIA 19.038 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.143 19.083 29.177 ;
      VIA 19.038 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.603 19.083 28.637 ;
      VIA 19.038 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.063 19.083 28.097 ;
      VIA 19.038 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 27.523 19.083 27.557 ;
      VIA 19.038 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.983 19.083 27.017 ;
      VIA 19.038 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.443 19.083 26.477 ;
      VIA 19.038 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.903 19.083 25.937 ;
      VIA 19.038 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.363 19.083 25.397 ;
      VIA 19.038 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.823 19.083 24.857 ;
      VIA 19.038 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.283 19.083 24.317 ;
      VIA 19.038 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.743 19.083 23.777 ;
      VIA 19.038 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.203 19.083 23.237 ;
      VIA 19.038 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.663 19.083 22.697 ;
      VIA 19.038 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.123 19.083 22.157 ;
      VIA 19.038 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.583 19.083 21.617 ;
      VIA 19.038 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.043 19.083 21.077 ;
      VIA 19.038 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 20.503 19.083 20.537 ;
      VIA 19.038 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.963 19.083 19.997 ;
      VIA 19.038 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.423 19.083 19.457 ;
      VIA 19.038 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.883 19.083 18.917 ;
      VIA 19.038 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.343 19.083 18.377 ;
      VIA 19.038 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.803 19.083 17.837 ;
      VIA 19.038 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.263 19.083 17.297 ;
      VIA 19.038 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.723 19.083 16.757 ;
      VIA 19.038 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.183 19.083 16.217 ;
      VIA 19.038 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.643 19.083 15.677 ;
      VIA 19.038 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.103 19.083 15.137 ;
      VIA 19.038 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.563 19.083 14.597 ;
      VIA 19.038 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.023 19.083 14.057 ;
      VIA 19.038 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 13.483 19.083 13.517 ;
      VIA 19.038 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.943 19.083 12.977 ;
      VIA 19.038 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.403 19.083 12.437 ;
      VIA 19.038 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.863 19.083 11.897 ;
      VIA 19.038 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.323 19.083 11.357 ;
      VIA 19.038 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.783 19.083 10.817 ;
      VIA 19.038 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.243 19.083 10.277 ;
      VIA 19.038 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.703 19.083 9.737 ;
      VIA 19.038 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.163 19.083 9.197 ;
      VIA 19.038 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.623 19.083 8.657 ;
      VIA 19.038 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.083 19.083 8.117 ;
      VIA 19.038 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.543 19.083 7.577 ;
      VIA 19.038 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.003 19.083 7.037 ;
      VIA 19.038 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 6.463 19.083 6.497 ;
      VIA 19.038 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.923 19.083 5.957 ;
      VIA 19.038 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.383 19.083 5.417 ;
      VIA 19.038 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.843 19.083 4.877 ;
      VIA 19.038 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.303 19.083 4.337 ;
      VIA 19.038 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.763 19.083 3.797 ;
      VIA 19.038 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.223 19.083 3.257 ;
      VIA 19.038 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.683 19.083 2.717 ;
      VIA 19.038 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.143 19.083 2.177 ;
      VIA 19.038 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.603 19.083 1.637 ;
      VIA 19.038 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.063 19.083 1.097 ;
      VIA 19.038 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 57.763 13.179 57.797 ;
      VIA 13.134 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 57.223 13.179 57.257 ;
      VIA 13.134 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 56.683 13.179 56.717 ;
      VIA 13.134 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 56.143 13.179 56.177 ;
      VIA 13.134 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 55.603 13.179 55.637 ;
      VIA 13.134 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 55.063 13.179 55.097 ;
      VIA 13.134 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 54.523 13.179 54.557 ;
      VIA 13.134 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 53.983 13.179 54.017 ;
      VIA 13.134 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 53.443 13.179 53.477 ;
      VIA 13.134 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 52.903 13.179 52.937 ;
      VIA 13.134 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 52.363 13.179 52.397 ;
      VIA 13.134 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 51.823 13.179 51.857 ;
      VIA 13.134 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 51.283 13.179 51.317 ;
      VIA 13.134 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 50.743 13.179 50.777 ;
      VIA 13.134 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 50.203 13.179 50.237 ;
      VIA 13.134 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 49.663 13.179 49.697 ;
      VIA 13.134 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 49.123 13.179 49.157 ;
      VIA 13.134 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 48.583 13.179 48.617 ;
      VIA 13.134 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 48.043 13.179 48.077 ;
      VIA 13.134 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 47.503 13.179 47.537 ;
      VIA 13.134 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 46.963 13.179 46.997 ;
      VIA 13.134 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 46.423 13.179 46.457 ;
      VIA 13.134 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 45.883 13.179 45.917 ;
      VIA 13.134 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 45.343 13.179 45.377 ;
      VIA 13.134 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 44.803 13.179 44.837 ;
      VIA 13.134 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 44.263 13.179 44.297 ;
      VIA 13.134 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 43.723 13.179 43.757 ;
      VIA 13.134 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 43.183 13.179 43.217 ;
      VIA 13.134 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 42.643 13.179 42.677 ;
      VIA 13.134 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 42.103 13.179 42.137 ;
      VIA 13.134 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 41.563 13.179 41.597 ;
      VIA 13.134 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 41.023 13.179 41.057 ;
      VIA 13.134 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 40.483 13.179 40.517 ;
      VIA 13.134 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.943 13.179 39.977 ;
      VIA 13.134 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.403 13.179 39.437 ;
      VIA 13.134 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.863 13.179 38.897 ;
      VIA 13.134 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.323 13.179 38.357 ;
      VIA 13.134 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.783 13.179 37.817 ;
      VIA 13.134 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.243 13.179 37.277 ;
      VIA 13.134 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.703 13.179 36.737 ;
      VIA 13.134 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.163 13.179 36.197 ;
      VIA 13.134 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.623 13.179 35.657 ;
      VIA 13.134 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.083 13.179 35.117 ;
      VIA 13.134 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.543 13.179 34.577 ;
      VIA 13.134 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.003 13.179 34.037 ;
      VIA 13.134 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 33.463 13.179 33.497 ;
      VIA 13.134 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.923 13.179 32.957 ;
      VIA 13.134 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.383 13.179 32.417 ;
      VIA 13.134 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.843 13.179 31.877 ;
      VIA 13.134 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.303 13.179 31.337 ;
      VIA 13.134 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.763 13.179 30.797 ;
      VIA 13.134 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.223 13.179 30.257 ;
      VIA 13.134 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.683 13.179 29.717 ;
      VIA 13.134 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.143 13.179 29.177 ;
      VIA 13.134 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.603 13.179 28.637 ;
      VIA 13.134 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.063 13.179 28.097 ;
      VIA 13.134 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 27.523 13.179 27.557 ;
      VIA 13.134 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.983 13.179 27.017 ;
      VIA 13.134 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.443 13.179 26.477 ;
      VIA 13.134 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.903 13.179 25.937 ;
      VIA 13.134 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.363 13.179 25.397 ;
      VIA 13.134 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.823 13.179 24.857 ;
      VIA 13.134 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.283 13.179 24.317 ;
      VIA 13.134 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.743 13.179 23.777 ;
      VIA 13.134 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.203 13.179 23.237 ;
      VIA 13.134 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.663 13.179 22.697 ;
      VIA 13.134 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.123 13.179 22.157 ;
      VIA 13.134 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.583 13.179 21.617 ;
      VIA 13.134 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.043 13.179 21.077 ;
      VIA 13.134 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 20.503 13.179 20.537 ;
      VIA 13.134 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.963 13.179 19.997 ;
      VIA 13.134 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.423 13.179 19.457 ;
      VIA 13.134 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.883 13.179 18.917 ;
      VIA 13.134 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.343 13.179 18.377 ;
      VIA 13.134 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.803 13.179 17.837 ;
      VIA 13.134 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.263 13.179 17.297 ;
      VIA 13.134 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.723 13.179 16.757 ;
      VIA 13.134 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.183 13.179 16.217 ;
      VIA 13.134 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.643 13.179 15.677 ;
      VIA 13.134 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.103 13.179 15.137 ;
      VIA 13.134 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.563 13.179 14.597 ;
      VIA 13.134 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.023 13.179 14.057 ;
      VIA 13.134 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 13.483 13.179 13.517 ;
      VIA 13.134 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.943 13.179 12.977 ;
      VIA 13.134 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.403 13.179 12.437 ;
      VIA 13.134 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.863 13.179 11.897 ;
      VIA 13.134 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.323 13.179 11.357 ;
      VIA 13.134 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.783 13.179 10.817 ;
      VIA 13.134 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.243 13.179 10.277 ;
      VIA 13.134 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.703 13.179 9.737 ;
      VIA 13.134 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.163 13.179 9.197 ;
      VIA 13.134 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.623 13.179 8.657 ;
      VIA 13.134 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.083 13.179 8.117 ;
      VIA 13.134 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.543 13.179 7.577 ;
      VIA 13.134 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.003 13.179 7.037 ;
      VIA 13.134 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 6.463 13.179 6.497 ;
      VIA 13.134 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.923 13.179 5.957 ;
      VIA 13.134 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.383 13.179 5.417 ;
      VIA 13.134 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.843 13.179 4.877 ;
      VIA 13.134 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.303 13.179 4.337 ;
      VIA 13.134 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.763 13.179 3.797 ;
      VIA 13.134 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.223 13.179 3.257 ;
      VIA 13.134 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.683 13.179 2.717 ;
      VIA 13.134 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.143 13.179 2.177 ;
      VIA 13.134 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.603 13.179 1.637 ;
      VIA 13.134 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.063 13.179 1.097 ;
      VIA 13.134 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 57.763 7.275 57.797 ;
      VIA 7.23 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 57.223 7.275 57.257 ;
      VIA 7.23 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 56.683 7.275 56.717 ;
      VIA 7.23 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 56.143 7.275 56.177 ;
      VIA 7.23 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 55.603 7.275 55.637 ;
      VIA 7.23 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 55.063 7.275 55.097 ;
      VIA 7.23 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 54.523 7.275 54.557 ;
      VIA 7.23 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 53.983 7.275 54.017 ;
      VIA 7.23 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 53.443 7.275 53.477 ;
      VIA 7.23 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 52.903 7.275 52.937 ;
      VIA 7.23 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 52.363 7.275 52.397 ;
      VIA 7.23 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 51.823 7.275 51.857 ;
      VIA 7.23 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 51.283 7.275 51.317 ;
      VIA 7.23 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 50.743 7.275 50.777 ;
      VIA 7.23 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 50.203 7.275 50.237 ;
      VIA 7.23 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 49.663 7.275 49.697 ;
      VIA 7.23 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 49.123 7.275 49.157 ;
      VIA 7.23 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 48.583 7.275 48.617 ;
      VIA 7.23 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 48.043 7.275 48.077 ;
      VIA 7.23 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 47.503 7.275 47.537 ;
      VIA 7.23 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 46.963 7.275 46.997 ;
      VIA 7.23 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 46.423 7.275 46.457 ;
      VIA 7.23 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 45.883 7.275 45.917 ;
      VIA 7.23 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 45.343 7.275 45.377 ;
      VIA 7.23 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 44.803 7.275 44.837 ;
      VIA 7.23 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 44.263 7.275 44.297 ;
      VIA 7.23 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 43.723 7.275 43.757 ;
      VIA 7.23 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 43.183 7.275 43.217 ;
      VIA 7.23 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 42.643 7.275 42.677 ;
      VIA 7.23 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 42.103 7.275 42.137 ;
      VIA 7.23 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 41.563 7.275 41.597 ;
      VIA 7.23 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 41.023 7.275 41.057 ;
      VIA 7.23 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 40.483 7.275 40.517 ;
      VIA 7.23 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.943 7.275 39.977 ;
      VIA 7.23 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.403 7.275 39.437 ;
      VIA 7.23 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.863 7.275 38.897 ;
      VIA 7.23 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.323 7.275 38.357 ;
      VIA 7.23 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.783 7.275 37.817 ;
      VIA 7.23 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.243 7.275 37.277 ;
      VIA 7.23 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.703 7.275 36.737 ;
      VIA 7.23 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.163 7.275 36.197 ;
      VIA 7.23 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.623 7.275 35.657 ;
      VIA 7.23 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.083 7.275 35.117 ;
      VIA 7.23 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.543 7.275 34.577 ;
      VIA 7.23 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.003 7.275 34.037 ;
      VIA 7.23 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 33.463 7.275 33.497 ;
      VIA 7.23 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.923 7.275 32.957 ;
      VIA 7.23 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.383 7.275 32.417 ;
      VIA 7.23 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.843 7.275 31.877 ;
      VIA 7.23 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.303 7.275 31.337 ;
      VIA 7.23 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.763 7.275 30.797 ;
      VIA 7.23 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.223 7.275 30.257 ;
      VIA 7.23 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.683 7.275 29.717 ;
      VIA 7.23 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.143 7.275 29.177 ;
      VIA 7.23 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.603 7.275 28.637 ;
      VIA 7.23 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.063 7.275 28.097 ;
      VIA 7.23 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 27.523 7.275 27.557 ;
      VIA 7.23 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.983 7.275 27.017 ;
      VIA 7.23 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.443 7.275 26.477 ;
      VIA 7.23 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.903 7.275 25.937 ;
      VIA 7.23 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.363 7.275 25.397 ;
      VIA 7.23 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.823 7.275 24.857 ;
      VIA 7.23 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.283 7.275 24.317 ;
      VIA 7.23 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.743 7.275 23.777 ;
      VIA 7.23 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.203 7.275 23.237 ;
      VIA 7.23 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.663 7.275 22.697 ;
      VIA 7.23 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.123 7.275 22.157 ;
      VIA 7.23 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.583 7.275 21.617 ;
      VIA 7.23 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.043 7.275 21.077 ;
      VIA 7.23 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 20.503 7.275 20.537 ;
      VIA 7.23 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.963 7.275 19.997 ;
      VIA 7.23 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.423 7.275 19.457 ;
      VIA 7.23 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.883 7.275 18.917 ;
      VIA 7.23 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.343 7.275 18.377 ;
      VIA 7.23 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.803 7.275 17.837 ;
      VIA 7.23 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.263 7.275 17.297 ;
      VIA 7.23 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.723 7.275 16.757 ;
      VIA 7.23 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.183 7.275 16.217 ;
      VIA 7.23 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.643 7.275 15.677 ;
      VIA 7.23 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.103 7.275 15.137 ;
      VIA 7.23 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.563 7.275 14.597 ;
      VIA 7.23 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.023 7.275 14.057 ;
      VIA 7.23 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 13.483 7.275 13.517 ;
      VIA 7.23 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.943 7.275 12.977 ;
      VIA 7.23 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.403 7.275 12.437 ;
      VIA 7.23 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.863 7.275 11.897 ;
      VIA 7.23 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.323 7.275 11.357 ;
      VIA 7.23 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.783 7.275 10.817 ;
      VIA 7.23 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.243 7.275 10.277 ;
      VIA 7.23 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.703 7.275 9.737 ;
      VIA 7.23 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.163 7.275 9.197 ;
      VIA 7.23 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.623 7.275 8.657 ;
      VIA 7.23 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.083 7.275 8.117 ;
      VIA 7.23 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.543 7.275 7.577 ;
      VIA 7.23 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.003 7.275 7.037 ;
      VIA 7.23 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 6.463 7.275 6.497 ;
      VIA 7.23 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.923 7.275 5.957 ;
      VIA 7.23 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.383 7.275 5.417 ;
      VIA 7.23 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.843 7.275 4.877 ;
      VIA 7.23 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.303 7.275 4.337 ;
      VIA 7.23 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.763 7.275 3.797 ;
      VIA 7.23 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.223 7.275 3.257 ;
      VIA 7.23 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.683 7.275 2.717 ;
      VIA 7.23 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.143 7.275 2.177 ;
      VIA 7.23 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.603 7.275 1.637 ;
      VIA 7.23 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.063 7.275 1.097 ;
      VIA 7.23 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 57.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 57.763 1.371 57.797 ;
      VIA 1.326 57.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 57.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 57.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 57.223 1.371 57.257 ;
      VIA 1.326 57.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 57.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 56.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 56.683 1.371 56.717 ;
      VIA 1.326 56.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 56.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 56.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 56.143 1.371 56.177 ;
      VIA 1.326 56.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 56.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 55.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 55.603 1.371 55.637 ;
      VIA 1.326 55.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 55.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 55.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 55.063 1.371 55.097 ;
      VIA 1.326 55.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 55.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 54.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 54.523 1.371 54.557 ;
      VIA 1.326 54.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 54.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 53.983 1.371 54.017 ;
      VIA 1.326 54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 53.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 53.443 1.371 53.477 ;
      VIA 1.326 53.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 53.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 52.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 52.903 1.371 52.937 ;
      VIA 1.326 52.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 52.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 52.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 52.363 1.371 52.397 ;
      VIA 1.326 52.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 52.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 51.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 51.823 1.371 51.857 ;
      VIA 1.326 51.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 51.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 51.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 51.283 1.371 51.317 ;
      VIA 1.326 51.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 51.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 50.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 50.743 1.371 50.777 ;
      VIA 1.326 50.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 50.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 50.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 50.203 1.371 50.237 ;
      VIA 1.326 50.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 50.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 49.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 49.663 1.371 49.697 ;
      VIA 1.326 49.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 49.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 49.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 49.123 1.371 49.157 ;
      VIA 1.326 49.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 49.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 48.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 48.583 1.371 48.617 ;
      VIA 1.326 48.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 48.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 48.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 48.043 1.371 48.077 ;
      VIA 1.326 48.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 48.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 47.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 47.503 1.371 47.537 ;
      VIA 1.326 47.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 47.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 46.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 46.963 1.371 46.997 ;
      VIA 1.326 46.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 46.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 46.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 46.423 1.371 46.457 ;
      VIA 1.326 46.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 46.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 45.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 45.883 1.371 45.917 ;
      VIA 1.326 45.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 45.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 45.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 45.343 1.371 45.377 ;
      VIA 1.326 45.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 45.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 44.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 44.803 1.371 44.837 ;
      VIA 1.326 44.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 44.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 44.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 44.263 1.371 44.297 ;
      VIA 1.326 44.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 44.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 43.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 43.723 1.371 43.757 ;
      VIA 1.326 43.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 43.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 43.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 43.183 1.371 43.217 ;
      VIA 1.326 43.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 43.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 42.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 42.643 1.371 42.677 ;
      VIA 1.326 42.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 42.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 42.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 42.103 1.371 42.137 ;
      VIA 1.326 42.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 42.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 41.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 41.563 1.371 41.597 ;
      VIA 1.326 41.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 41.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 41.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 41.023 1.371 41.057 ;
      VIA 1.326 41.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 41.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 40.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 40.483 1.371 40.517 ;
      VIA 1.326 40.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 40.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.943 1.371 39.977 ;
      VIA 1.326 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.403 1.371 39.437 ;
      VIA 1.326 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.863 1.371 38.897 ;
      VIA 1.326 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.323 1.371 38.357 ;
      VIA 1.326 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.783 1.371 37.817 ;
      VIA 1.326 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.243 1.371 37.277 ;
      VIA 1.326 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.703 1.371 36.737 ;
      VIA 1.326 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.163 1.371 36.197 ;
      VIA 1.326 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.623 1.371 35.657 ;
      VIA 1.326 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.083 1.371 35.117 ;
      VIA 1.326 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.543 1.371 34.577 ;
      VIA 1.326 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.003 1.371 34.037 ;
      VIA 1.326 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 33.463 1.371 33.497 ;
      VIA 1.326 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.923 1.371 32.957 ;
      VIA 1.326 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.383 1.371 32.417 ;
      VIA 1.326 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.843 1.371 31.877 ;
      VIA 1.326 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.303 1.371 31.337 ;
      VIA 1.326 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.763 1.371 30.797 ;
      VIA 1.326 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.223 1.371 30.257 ;
      VIA 1.326 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.683 1.371 29.717 ;
      VIA 1.326 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.143 1.371 29.177 ;
      VIA 1.326 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.603 1.371 28.637 ;
      VIA 1.326 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.063 1.371 28.097 ;
      VIA 1.326 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 27.523 1.371 27.557 ;
      VIA 1.326 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.983 1.371 27.017 ;
      VIA 1.326 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.443 1.371 26.477 ;
      VIA 1.326 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.903 1.371 25.937 ;
      VIA 1.326 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.363 1.371 25.397 ;
      VIA 1.326 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.823 1.371 24.857 ;
      VIA 1.326 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.283 1.371 24.317 ;
      VIA 1.326 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.743 1.371 23.777 ;
      VIA 1.326 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.203 1.371 23.237 ;
      VIA 1.326 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.663 1.371 22.697 ;
      VIA 1.326 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.123 1.371 22.157 ;
      VIA 1.326 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.583 1.371 21.617 ;
      VIA 1.326 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.043 1.371 21.077 ;
      VIA 1.326 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 20.503 1.371 20.537 ;
      VIA 1.326 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.963 1.371 19.997 ;
      VIA 1.326 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.423 1.371 19.457 ;
      VIA 1.326 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.883 1.371 18.917 ;
      VIA 1.326 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.343 1.371 18.377 ;
      VIA 1.326 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.803 1.371 17.837 ;
      VIA 1.326 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.263 1.371 17.297 ;
      VIA 1.326 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.723 1.371 16.757 ;
      VIA 1.326 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.183 1.371 16.217 ;
      VIA 1.326 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.643 1.371 15.677 ;
      VIA 1.326 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.103 1.371 15.137 ;
      VIA 1.326 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.563 1.371 14.597 ;
      VIA 1.326 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.023 1.371 14.057 ;
      VIA 1.326 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 13.483 1.371 13.517 ;
      VIA 1.326 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.943 1.371 12.977 ;
      VIA 1.326 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.403 1.371 12.437 ;
      VIA 1.326 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.863 1.371 11.897 ;
      VIA 1.326 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.323 1.371 11.357 ;
      VIA 1.326 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.783 1.371 10.817 ;
      VIA 1.326 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.243 1.371 10.277 ;
      VIA 1.326 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.703 1.371 9.737 ;
      VIA 1.326 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.163 1.371 9.197 ;
      VIA 1.326 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.623 1.371 8.657 ;
      VIA 1.326 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.083 1.371 8.117 ;
      VIA 1.326 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.543 1.371 7.577 ;
      VIA 1.326 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.003 1.371 7.037 ;
      VIA 1.326 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 6.463 1.371 6.497 ;
      VIA 1.326 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.923 1.371 5.957 ;
      VIA 1.326 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.383 1.371 5.417 ;
      VIA 1.326 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 29.565 57.78 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 57.24 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 56.7 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 56.16 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 55.62 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 55.08 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 54.54 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 54 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 53.46 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 52.92 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 52.38 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 51.84 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 51.3 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 50.76 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 50.22 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 49.68 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 49.14 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 48.6 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 48.06 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 47.52 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 46.98 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 46.44 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 45.9 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 45.36 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 44.82 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 44.28 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 43.74 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 43.2 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 42.66 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 42.12 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 41.58 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 41.04 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 40.5 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 39.96 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 39.42 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 38.88 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 38.34 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 37.8 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 37.26 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 36.72 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 36.18 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 35.64 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 35.1 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 34.56 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 34.02 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 33.48 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 32.94 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 32.4 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 31.86 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 31.32 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 30.78 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 30.24 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 29.7 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 29.16 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 28.62 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 28.08 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 27.54 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 27 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 26.46 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 25.92 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 25.38 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 24.84 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 24.3 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 23.76 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 23.22 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 22.68 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 22.14 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 21.6 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 21.06 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 20.52 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 19.98 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 19.44 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 18.9 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 18.36 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 17.82 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 17.28 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 16.74 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 16.2 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 15.66 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 15.12 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 14.58 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 14.04 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 13.5 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 12.96 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 12.42 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 11.88 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 11.34 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 10.8 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 10.26 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 9.72 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 9.18 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 8.64 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 8.1 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 7.56 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 7.02 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 6.48 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 5.94 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 5.4 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 4.86 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 4.32 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 3.78 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 3.24 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 2.7 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 2.16 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 1.62 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
      VIA 29.565 1.08 run_benchmark_via1_2_57078_18_1_1585_36_36 ;
    END
  END VSS
  PIN M_DataRdy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.672 0 0.696 0.084 ;
    END
  END M_DataRdy[0]
  PIN M_DataRdy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.768 0 0.792 0.084 ;
    END
  END M_DataRdy[1]
  PIN M_Rdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.232 0 23.256 0.084 ;
    END
  END M_Rdata_ram[0]
  PIN M_Rdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.88 0 26.904 0.084 ;
    END
  END M_Rdata_ram[10]
  PIN M_Rdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.408 0 21.432 0.084 ;
    END
  END M_Rdata_ram[11]
  PIN M_Rdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.976 0 27 0.084 ;
    END
  END M_Rdata_ram[12]
  PIN M_Rdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.416 0 28.44 0.084 ;
    END
  END M_Rdata_ram[13]
  PIN M_Rdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.648 0 27.672 0.084 ;
    END
  END M_Rdata_ram[14]
  PIN M_Rdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.448 0 20.472 0.084 ;
    END
  END M_Rdata_ram[15]
  PIN M_Rdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.928 0 20.952 0.084 ;
    END
  END M_Rdata_ram[16]
  PIN M_Rdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.64 0 20.664 0.084 ;
    END
  END M_Rdata_ram[17]
  PIN M_Rdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.872 0 19.896 0.084 ;
    END
  END M_Rdata_ram[18]
  PIN M_Rdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.704 0 28.728 0.084 ;
    END
  END M_Rdata_ram[19]
  PIN M_Rdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 0 21.72 0.084 ;
    END
  END M_Rdata_ram[1]
  PIN M_Rdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.064 0 20.088 0.084 ;
    END
  END M_Rdata_ram[20]
  PIN M_Rdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.904 0 35.928 0.084 ;
    END
  END M_Rdata_ram[21]
  PIN M_Rdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.808 0 35.832 0.084 ;
    END
  END M_Rdata_ram[22]
  PIN M_Rdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.712 0 35.736 0.084 ;
    END
  END M_Rdata_ram[23]
  PIN M_Rdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.616 0 35.64 0.084 ;
    END
  END M_Rdata_ram[24]
  PIN M_Rdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.832 0 32.856 0.084 ;
    END
  END M_Rdata_ram[25]
  PIN M_Rdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.584 0 31.608 0.084 ;
    END
  END M_Rdata_ram[26]
  PIN M_Rdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.776 0 31.8 0.084 ;
    END
  END M_Rdata_ram[27]
  PIN M_Rdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.816 0 30.84 0.084 ;
    END
  END M_Rdata_ram[28]
  PIN M_Rdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.856 0 29.88 0.084 ;
    END
  END M_Rdata_ram[29]
  PIN M_Rdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.56 0 22.584 0.084 ;
    END
  END M_Rdata_ram[2]
  PIN M_Rdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.144 0 30.168 0.084 ;
    END
  END M_Rdata_ram[30]
  PIN M_Rdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.032 0 28.056 0.084 ;
    END
  END M_Rdata_ram[31]
  PIN M_Rdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.728 0 25.752 0.084 ;
    END
  END M_Rdata_ram[32]
  PIN M_Rdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.328 0 23.352 0.084 ;
    END
  END M_Rdata_ram[33]
  PIN M_Rdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.712 0 23.736 0.084 ;
    END
  END M_Rdata_ram[34]
  PIN M_Rdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.136 0 23.16 0.084 ;
    END
  END M_Rdata_ram[35]
  PIN M_Rdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.848 0 22.872 0.084 ;
    END
  END M_Rdata_ram[36]
  PIN M_Rdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.632 0 25.656 0.084 ;
    END
  END M_Rdata_ram[37]
  PIN M_Rdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.152 0 25.176 0.084 ;
    END
  END M_Rdata_ram[38]
  PIN M_Rdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.672 0 24.696 0.084 ;
    END
  END M_Rdata_ram[39]
  PIN M_Rdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.656 0 22.68 0.084 ;
    END
  END M_Rdata_ram[3]
  PIN M_Rdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.184 0 29.208 0.084 ;
    END
  END M_Rdata_ram[40]
  PIN M_Rdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.376 0 29.4 0.084 ;
    END
  END M_Rdata_ram[41]
  PIN M_Rdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.28 0 29.304 0.084 ;
    END
  END M_Rdata_ram[42]
  PIN M_Rdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.72 0 30.744 0.084 ;
    END
  END M_Rdata_ram[43]
  PIN M_Rdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.912 0 30.936 0.084 ;
    END
  END M_Rdata_ram[44]
  PIN M_Rdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.8 0 28.824 0.084 ;
    END
  END M_Rdata_ram[45]
  PIN M_Rdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.064 0 32.088 0.084 ;
    END
  END M_Rdata_ram[46]
  PIN M_Rdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.576 0 24.6 0.084 ;
    END
  END M_Rdata_ram[47]
  PIN M_Rdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.888 0 33.912 0.084 ;
    END
  END M_Rdata_ram[48]
  PIN M_Rdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.36 0 27.384 0.084 ;
    END
  END M_Rdata_ram[49]
  PIN M_Rdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.52 0 23.544 0.084 ;
    END
  END M_Rdata_ram[4]
  PIN M_Rdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.52 0 35.544 0.084 ;
    END
  END M_Rdata_ram[50]
  PIN M_Rdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.176 0 34.2 0.084 ;
    END
  END M_Rdata_ram[51]
  PIN M_Rdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.272 0 34.296 0.084 ;
    END
  END M_Rdata_ram[52]
  PIN M_Rdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.656 0 34.68 0.084 ;
    END
  END M_Rdata_ram[53]
  PIN M_Rdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.04 0 35.064 0.084 ;
    END
  END M_Rdata_ram[54]
  PIN M_Rdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.424 0 35.448 0.084 ;
    END
  END M_Rdata_ram[55]
  PIN M_Rdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.328 0 35.352 0.084 ;
    END
  END M_Rdata_ram[56]
  PIN M_Rdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.968 0 31.992 0.084 ;
    END
  END M_Rdata_ram[57]
  PIN M_Rdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.496 0 26.52 0.084 ;
    END
  END M_Rdata_ram[58]
  PIN M_Rdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.736 0 32.76 0.084 ;
    END
  END M_Rdata_ram[59]
  PIN M_Rdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.12 0 21.144 0.084 ;
    END
  END M_Rdata_ram[5]
  PIN M_Rdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.76 0 29.784 0.084 ;
    END
  END M_Rdata_ram[60]
  PIN M_Rdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.048 0 30.072 0.084 ;
    END
  END M_Rdata_ram[61]
  PIN M_Rdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.432 0 30.456 0.084 ;
    END
  END M_Rdata_ram[62]
  PIN M_Rdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.176 0 22.2 0.084 ;
    END
  END M_Rdata_ram[63]
  PIN M_Rdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.288 0 24.312 0.084 ;
    END
  END M_Rdata_ram[6]
  PIN M_Rdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.4 0 26.424 0.084 ;
    END
  END M_Rdata_ram[7]
  PIN M_Rdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.072 0 27.096 0.084 ;
    END
  END M_Rdata_ram[8]
  PIN M_Rdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.736 0 20.76 0.084 ;
    END
  END M_Rdata_ram[9]
  PIN Min_Wdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.592 0 26.616 0.084 ;
    END
  END Min_Wdata_ram[0]
  PIN Min_Wdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.24 0 30.264 0.084 ;
    END
  END Min_Wdata_ram[10]
  PIN Min_Wdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.504 0 33.528 0.084 ;
    END
  END Min_Wdata_ram[11]
  PIN Min_Wdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.544 0 32.568 0.084 ;
    END
  END Min_Wdata_ram[12]
  PIN Min_Wdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.408 0 33.432 0.084 ;
    END
  END Min_Wdata_ram[13]
  PIN Min_Wdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.944 0 34.968 0.084 ;
    END
  END Min_Wdata_ram[14]
  PIN Min_Wdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.48 0 36.504 0.084 ;
    END
  END Min_Wdata_ram[15]
  PIN Min_Wdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.76 0 41.784 0.084 ;
    END
  END Min_Wdata_ram[16]
  PIN Min_Wdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.88 0 38.904 0.084 ;
    END
  END Min_Wdata_ram[17]
  PIN Min_Wdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.28 0 41.304 0.084 ;
    END
  END Min_Wdata_ram[18]
  PIN Min_Wdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.184 0 41.208 0.084 ;
    END
  END Min_Wdata_ram[19]
  PIN Min_Wdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.48 0 24.504 0.084 ;
    END
  END Min_Wdata_ram[1]
  PIN Min_Wdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.936 0 39.96 0.084 ;
    END
  END Min_Wdata_ram[20]
  PIN Min_Wdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.664 0 41.688 0.084 ;
    END
  END Min_Wdata_ram[21]
  PIN Min_Wdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.896 0 40.92 0.084 ;
    END
  END Min_Wdata_ram[22]
  PIN Min_Wdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.512 0 40.536 0.084 ;
    END
  END Min_Wdata_ram[23]
  PIN Min_Wdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.648 0 39.672 0.084 ;
    END
  END Min_Wdata_ram[24]
  PIN Min_Wdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.976 0 39 0.084 ;
    END
  END Min_Wdata_ram[25]
  PIN Min_Wdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.112 0 38.136 0.084 ;
    END
  END Min_Wdata_ram[26]
  PIN Min_Wdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.192 0 36.216 0.084 ;
    END
  END Min_Wdata_ram[27]
  PIN Min_Wdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.464 0 34.488 0.084 ;
    END
  END Min_Wdata_ram[28]
  PIN Min_Wdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.336 0 30.36 0.084 ;
    END
  END Min_Wdata_ram[29]
  PIN Min_Wdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.272 0 22.296 0.084 ;
    END
  END Min_Wdata_ram[2]
  PIN Min_Wdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.64 0 32.664 0.084 ;
    END
  END Min_Wdata_ram[30]
  PIN Min_Wdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.128 0 28.152 0.084 ;
    END
  END Min_Wdata_ram[31]
  PIN Min_Wdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.6 0 21.624 0.084 ;
    END
  END Min_Wdata_ram[32]
  PIN Min_Wdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.168 0 27.192 0.084 ;
    END
  END Min_Wdata_ram[33]
  PIN Min_Wdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.936 0 27.96 0.084 ;
    END
  END Min_Wdata_ram[34]
  PIN Min_Wdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.344 0 25.368 0.084 ;
    END
  END Min_Wdata_ram[35]
  PIN Min_Wdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.536 0 25.56 0.084 ;
    END
  END Min_Wdata_ram[36]
  PIN Min_Wdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.264 0 27.288 0.084 ;
    END
  END Min_Wdata_ram[37]
  PIN Min_Wdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.04 0 23.064 0.084 ;
    END
  END Min_Wdata_ram[38]
  PIN Min_Wdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.896 0 28.92 0.084 ;
    END
  END Min_Wdata_ram[39]
  PIN Min_Wdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.944 0 22.968 0.084 ;
    END
  END Min_Wdata_ram[3]
  PIN Min_Wdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.2 0 31.224 0.084 ;
    END
  END Min_Wdata_ram[40]
  PIN Min_Wdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.488 0 31.512 0.084 ;
    END
  END Min_Wdata_ram[41]
  PIN Min_Wdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.664 0 29.688 0.084 ;
    END
  END Min_Wdata_ram[42]
  PIN Min_Wdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.216 0 33.24 0.084 ;
    END
  END Min_Wdata_ram[43]
  PIN Min_Wdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.256 0 32.28 0.084 ;
    END
  END Min_Wdata_ram[44]
  PIN Min_Wdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.696 0 33.72 0.084 ;
    END
  END Min_Wdata_ram[45]
  PIN Min_Wdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.848 0 34.872 0.084 ;
    END
  END Min_Wdata_ram[46]
  PIN Min_Wdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.576 0 36.6 0.084 ;
    END
  END Min_Wdata_ram[47]
  PIN Min_Wdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.864 0 36.888 0.084 ;
    END
  END Min_Wdata_ram[48]
  PIN Min_Wdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.96 0 36.984 0.084 ;
    END
  END Min_Wdata_ram[49]
  PIN Min_Wdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.752 0 22.776 0.084 ;
    END
  END Min_Wdata_ram[4]
  PIN Min_Wdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.728 0 37.752 0.084 ;
    END
  END Min_Wdata_ram[50]
  PIN Min_Wdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.44 0 37.464 0.084 ;
    END
  END Min_Wdata_ram[51]
  PIN Min_Wdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.056 0 37.08 0.084 ;
    END
  END Min_Wdata_ram[52]
  PIN Min_Wdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.152 0 37.176 0.084 ;
    END
  END Min_Wdata_ram[53]
  PIN Min_Wdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.248 0 37.272 0.084 ;
    END
  END Min_Wdata_ram[54]
  PIN Min_Wdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.824 0 37.848 0.084 ;
    END
  END Min_Wdata_ram[55]
  PIN Min_Wdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.536 0 37.56 0.084 ;
    END
  END Min_Wdata_ram[56]
  PIN Min_Wdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.496 0 38.52 0.084 ;
    END
  END Min_Wdata_ram[57]
  PIN Min_Wdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36 0 36.024 0.084 ;
    END
  END Min_Wdata_ram[58]
  PIN Min_Wdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.368 0 34.392 0.084 ;
    END
  END Min_Wdata_ram[59]
  PIN Min_Wdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24 0 24.024 0.084 ;
    END
  END Min_Wdata_ram[5]
  PIN Min_Wdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.792 0 33.816 0.084 ;
    END
  END Min_Wdata_ram[60]
  PIN Min_Wdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.008 0 31.032 0.084 ;
    END
  END Min_Wdata_ram[61]
  PIN Min_Wdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.352 0 32.376 0.084 ;
    END
  END Min_Wdata_ram[62]
  PIN Min_Wdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.472 0 29.496 0.084 ;
    END
  END Min_Wdata_ram[63]
  PIN Min_Wdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.808 0 23.832 0.084 ;
    END
  END Min_Wdata_ram[6]
  PIN Min_Wdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.552 0 27.576 0.084 ;
    END
  END Min_Wdata_ram[7]
  PIN Min_Wdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.392 0 31.416 0.084 ;
    END
  END Min_Wdata_ram[8]
  PIN Min_Wdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.312 0 33.336 0.084 ;
    END
  END Min_Wdata_ram[9]
  PIN Min_addr_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.224 0 28.248 0.084 ;
    END
  END Min_addr_ram[0]
  PIN Min_addr_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.56 0.084 22.584 ;
    END
  END Min_addr_ram[10]
  PIN Min_addr_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.888 0 21.912 0.084 ;
    END
  END Min_addr_ram[11]
  PIN Min_addr_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.096 0 24.12 0.084 ;
    END
  END Min_addr_ram[12]
  PIN Min_addr_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.544 0 20.568 0.084 ;
    END
  END Min_addr_ram[13]
  PIN Min_addr_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.08 0 22.104 0.084 ;
    END
  END Min_addr_ram[14]
  PIN Min_addr_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.44 0 25.464 0.084 ;
    END
  END Min_addr_ram[15]
  PIN Min_addr_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.832 0 20.856 0.084 ;
    END
  END Min_addr_ram[16]
  PIN Min_addr_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.864 0 24.888 0.084 ;
    END
  END Min_addr_ram[17]
  PIN Min_addr_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.792 0 21.816 0.084 ;
    END
  END Min_addr_ram[18]
  PIN Min_addr_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.024 0 21.048 0.084 ;
    END
  END Min_addr_ram[19]
  PIN Min_addr_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.16 0 20.184 0.084 ;
    END
  END Min_addr_ram[1]
  PIN Min_addr_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.456 0 27.48 0.084 ;
    END
  END Min_addr_ram[20]
  PIN Min_addr_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.256 0 20.28 0.084 ;
    END
  END Min_addr_ram[21]
  PIN Min_addr_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.512 0 28.536 0.084 ;
    END
  END Min_addr_ram[22]
  PIN Min_addr_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.336 59.037 30.36 59.121 ;
    END
  END Min_addr_ram[23]
  PIN Min_addr_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.24 59.037 30.264 59.121 ;
    END
  END Min_addr_ram[24]
  PIN Min_addr_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.32 59.037 28.344 59.121 ;
    END
  END Min_addr_ram[25]
  PIN Min_addr_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.776 59.037 31.8 59.121 ;
    END
  END Min_addr_ram[26]
  PIN Min_addr_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.008 59.037 31.032 59.121 ;
    END
  END Min_addr_ram[27]
  PIN Min_addr_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.104 59.037 31.128 59.121 ;
    END
  END Min_addr_ram[28]
  PIN Min_addr_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.528 59.037 30.552 59.121 ;
    END
  END Min_addr_ram[29]
  PIN Min_addr_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.464 0 22.488 0.084 ;
    END
  END Min_addr_ram[2]
  PIN Min_addr_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.416 59.037 28.44 59.121 ;
    END
  END Min_addr_ram[30]
  PIN Min_addr_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.856 59.037 29.88 59.121 ;
    END
  END Min_addr_ram[31]
  PIN Min_addr_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.296 59.037 31.32 59.121 ;
    END
  END Min_addr_ram[32]
  PIN Min_addr_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.2 59.037 31.224 59.121 ;
    END
  END Min_addr_ram[33]
  PIN Min_addr_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.912 59.037 30.936 59.121 ;
    END
  END Min_addr_ram[34]
  PIN Min_addr_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.448 59.037 32.472 59.121 ;
    END
  END Min_addr_ram[35]
  PIN Min_addr_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.544 59.037 32.568 59.121 ;
    END
  END Min_addr_ram[36]
  PIN Min_addr_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.352 59.037 32.376 59.121 ;
    END
  END Min_addr_ram[37]
  PIN Min_addr_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.576 59.037 36.6 59.121 ;
    END
  END Min_addr_ram[38]
  PIN Min_addr_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.808 59.037 35.832 59.121 ;
    END
  END Min_addr_ram[39]
  PIN Min_addr_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.312 0 21.336 0.084 ;
    END
  END Min_addr_ram[3]
  PIN Min_addr_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.136 59.037 35.16 59.121 ;
    END
  END Min_addr_ram[40]
  PIN Min_addr_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.616 59.037 35.64 59.121 ;
    END
  END Min_addr_ram[41]
  PIN Min_addr_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.768 59.037 36.792 59.121 ;
    END
  END Min_addr_ram[42]
  PIN Min_addr_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.864 59.037 36.888 59.121 ;
    END
  END Min_addr_ram[43]
  PIN Min_addr_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.96 59.037 36.984 59.121 ;
    END
  END Min_addr_ram[44]
  PIN Min_addr_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.672 59.037 36.696 59.121 ;
    END
  END Min_addr_ram[45]
  PIN Min_addr_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.632 0.084 25.656 ;
    END
  END Min_addr_ram[4]
  PIN Min_addr_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.344 0.084 25.368 ;
    END
  END Min_addr_ram[5]
  PIN Min_addr_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.672 0.084 24.696 ;
    END
  END Min_addr_ram[6]
  PIN Min_addr_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.48 0.084 24.504 ;
    END
  END Min_addr_ram[7]
  PIN Min_addr_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.904 0.084 23.928 ;
    END
  END Min_addr_ram[8]
  PIN Min_addr_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.808 0.084 23.832 ;
    END
  END Min_addr_ram[9]
  PIN Min_data_ram_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.904 0 23.928 0.084 ;
    END
  END Min_data_ram_size[0]
  PIN Min_data_ram_size[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.704 59.037 28.728 59.121 ;
    END
  END Min_data_ram_size[10]
  PIN Min_data_ram_size[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.896 59.037 28.92 59.121 ;
    END
  END Min_data_ram_size[11]
  PIN Min_data_ram_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.352 0 20.376 0.084 ;
    END
  END Min_data_ram_size[1]
  PIN Min_data_ram_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.424 0 23.448 0.084 ;
    END
  END Min_data_ram_size[2]
  PIN Min_data_ram_size[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.824 0 25.848 0.084 ;
    END
  END Min_data_ram_size[3]
  PIN Min_data_ram_size[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.92 0 25.944 0.084 ;
    END
  END Min_data_ram_size[4]
  PIN Min_data_ram_size[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.84 0 27.864 0.084 ;
    END
  END Min_data_ram_size[5]
  PIN Min_data_ram_size[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.088 59.037 29.112 59.121 ;
    END
  END Min_data_ram_size[6]
  PIN Min_data_ram_size[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.512 59.037 28.536 59.121 ;
    END
  END Min_data_ram_size[7]
  PIN Min_data_ram_size[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.8 59.037 28.824 59.121 ;
    END
  END Min_data_ram_size[8]
  PIN Min_data_ram_size[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.184 59.037 29.208 59.121 ;
    END
  END Min_data_ram_size[9]
  PIN Min_oe_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.744 0 27.768 0.084 ;
    END
  END Min_oe_ram[0]
  PIN Min_oe_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.52 59.037 35.544 59.121 ;
    END
  END Min_oe_ram[1]
  PIN Min_we_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.968 0 19.992 0.084 ;
    END
  END Min_we_ram[0]
  PIN Min_we_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.608 59.037 28.632 59.121 ;
    END
  END Min_we_ram[1]
  PIN Mout_Wdata_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.384 0 24.408 0.084 ;
    END
  END Mout_Wdata_ram[0]
  PIN Mout_Wdata_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.624 0 30.648 0.084 ;
    END
  END Mout_Wdata_ram[10]
  PIN Mout_Wdata_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.616 0 23.64 0.084 ;
    END
  END Mout_Wdata_ram[11]
  PIN Mout_Wdata_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.872 0 31.896 0.084 ;
    END
  END Mout_Wdata_ram[12]
  PIN Mout_Wdata_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.984 0 34.008 0.084 ;
    END
  END Mout_Wdata_ram[13]
  PIN Mout_Wdata_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.232 0 35.256 0.084 ;
    END
  END Mout_Wdata_ram[14]
  PIN Mout_Wdata_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.288 0 36.312 0.084 ;
    END
  END Mout_Wdata_ram[15]
  PIN Mout_Wdata_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.744 0 39.768 0.084 ;
    END
  END Mout_Wdata_ram[16]
  PIN Mout_Wdata_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.568 0 41.592 0.084 ;
    END
  END Mout_Wdata_ram[17]
  PIN Mout_Wdata_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.608 0 40.632 0.084 ;
    END
  END Mout_Wdata_ram[18]
  PIN Mout_Wdata_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.088 0 41.112 0.084 ;
    END
  END Mout_Wdata_ram[19]
  PIN Mout_Wdata_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.056 0 25.08 0.084 ;
    END
  END Mout_Wdata_ram[1]
  PIN Mout_Wdata_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.416 0 40.44 0.084 ;
    END
  END Mout_Wdata_ram[20]
  PIN Mout_Wdata_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.032 0 40.056 0.084 ;
    END
  END Mout_Wdata_ram[21]
  PIN Mout_Wdata_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.224 0 40.248 0.084 ;
    END
  END Mout_Wdata_ram[22]
  PIN Mout_Wdata_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.128 0 40.152 0.084 ;
    END
  END Mout_Wdata_ram[23]
  PIN Mout_Wdata_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.376 0 41.4 0.084 ;
    END
  END Mout_Wdata_ram[24]
  PIN Mout_Wdata_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.32 0 40.344 0.084 ;
    END
  END Mout_Wdata_ram[25]
  PIN Mout_Wdata_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.304 0 38.328 0.084 ;
    END
  END Mout_Wdata_ram[26]
  PIN Mout_Wdata_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.384 0 36.408 0.084 ;
    END
  END Mout_Wdata_ram[27]
  PIN Mout_Wdata_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.752 0 34.776 0.084 ;
    END
  END Mout_Wdata_ram[28]
  PIN Mout_Wdata_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.528 0 30.552 0.084 ;
    END
  END Mout_Wdata_ram[29]
  PIN Mout_Wdata_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.768 0 24.792 0.084 ;
    END
  END Mout_Wdata_ram[2]
  PIN Mout_Wdata_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.928 0 32.952 0.084 ;
    END
  END Mout_Wdata_ram[30]
  PIN Mout_Wdata_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.088 0 29.112 0.084 ;
    END
  END Mout_Wdata_ram[31]
  PIN Mout_Wdata_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.504 0 21.528 0.084 ;
    END
  END Mout_Wdata_ram[32]
  PIN Mout_Wdata_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.208 0 26.232 0.084 ;
    END
  END Mout_Wdata_ram[33]
  PIN Mout_Wdata_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.608 0 28.632 0.084 ;
    END
  END Mout_Wdata_ram[34]
  PIN Mout_Wdata_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.304 0 26.328 0.084 ;
    END
  END Mout_Wdata_ram[35]
  PIN Mout_Wdata_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.688 0 26.712 0.084 ;
    END
  END Mout_Wdata_ram[36]
  PIN Mout_Wdata_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.784 0 26.808 0.084 ;
    END
  END Mout_Wdata_ram[37]
  PIN Mout_Wdata_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.992 0 29.016 0.084 ;
    END
  END Mout_Wdata_ram[38]
  PIN Mout_Wdata_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.368 0 22.392 0.084 ;
    END
  END Mout_Wdata_ram[39]
  PIN Mout_Wdata_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.96 0 24.984 0.084 ;
    END
  END Mout_Wdata_ram[3]
  PIN Mout_Wdata_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.296 0 31.32 0.084 ;
    END
  END Mout_Wdata_ram[40]
  PIN Mout_Wdata_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.12 0 33.144 0.084 ;
    END
  END Mout_Wdata_ram[41]
  PIN Mout_Wdata_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.952 0 29.976 0.084 ;
    END
  END Mout_Wdata_ram[42]
  PIN Mout_Wdata_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.024 0 33.048 0.084 ;
    END
  END Mout_Wdata_ram[43]
  PIN Mout_Wdata_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.448 0 32.472 0.084 ;
    END
  END Mout_Wdata_ram[44]
  PIN Mout_Wdata_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.016 0 26.04 0.084 ;
    END
  END Mout_Wdata_ram[45]
  PIN Mout_Wdata_ram[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.136 0 35.16 0.084 ;
    END
  END Mout_Wdata_ram[46]
  PIN Mout_Wdata_ram[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.672 0 36.696 0.084 ;
    END
  END Mout_Wdata_ram[47]
  PIN Mout_Wdata_ram[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.768 0 36.792 0.084 ;
    END
  END Mout_Wdata_ram[48]
  PIN Mout_Wdata_ram[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.688 0 38.712 0.084 ;
    END
  END Mout_Wdata_ram[49]
  PIN Mout_Wdata_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.216 0 21.24 0.084 ;
    END
  END Mout_Wdata_ram[4]
  PIN Mout_Wdata_ram[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.208 0 38.232 0.084 ;
    END
  END Mout_Wdata_ram[50]
  PIN Mout_Wdata_ram[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.632 0 37.656 0.084 ;
    END
  END Mout_Wdata_ram[51]
  PIN Mout_Wdata_ram[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.92 0 37.944 0.084 ;
    END
  END Mout_Wdata_ram[52]
  PIN Mout_Wdata_ram[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.344 0 37.368 0.084 ;
    END
  END Mout_Wdata_ram[53]
  PIN Mout_Wdata_ram[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.016 0 38.04 0.084 ;
    END
  END Mout_Wdata_ram[54]
  PIN Mout_Wdata_ram[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.784 0 38.808 0.084 ;
    END
  END Mout_Wdata_ram[55]
  PIN Mout_Wdata_ram[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.4 0 38.424 0.084 ;
    END
  END Mout_Wdata_ram[56]
  PIN Mout_Wdata_ram[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  38.592 0 38.616 0.084 ;
    END
  END Mout_Wdata_ram[57]
  PIN Mout_Wdata_ram[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.096 0 36.12 0.084 ;
    END
  END Mout_Wdata_ram[58]
  PIN Mout_Wdata_ram[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.56 0 34.584 0.084 ;
    END
  END Mout_Wdata_ram[59]
  PIN Mout_Wdata_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.192 0 24.216 0.084 ;
    END
  END Mout_Wdata_ram[5]
  PIN Mout_Wdata_ram[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  34.08 0 34.104 0.084 ;
    END
  END Mout_Wdata_ram[60]
  PIN Mout_Wdata_ram[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.104 0 31.128 0.084 ;
    END
  END Mout_Wdata_ram[61]
  PIN Mout_Wdata_ram[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.16 0 32.184 0.084 ;
    END
  END Mout_Wdata_ram[62]
  PIN Mout_Wdata_ram[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.568 0 29.592 0.084 ;
    END
  END Mout_Wdata_ram[63]
  PIN Mout_Wdata_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.112 0 26.136 0.084 ;
    END
  END Mout_Wdata_ram[6]
  PIN Mout_Wdata_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.32 0 28.344 0.084 ;
    END
  END Mout_Wdata_ram[7]
  PIN Mout_Wdata_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.68 0 31.704 0.084 ;
    END
  END Mout_Wdata_ram[8]
  PIN Mout_Wdata_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.6 0 33.624 0.084 ;
    END
  END Mout_Wdata_ram[9]
  PIN Mout_addr_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  25.248 0 25.272 0.084 ;
    END
  END Mout_addr_ram[0]
  PIN Mout_addr_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.368 0.084 22.392 ;
    END
  END Mout_addr_ram[10]
  PIN Mout_addr_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 0 22.008 0.084 ;
    END
  END Mout_addr_ram[11]
  PIN Mout_addr_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.696 0.084 21.72 ;
    END
  END Mout_addr_ram[12]
  PIN Mout_addr_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.928 0.084 20.952 ;
    END
  END Mout_addr_ram[13]
  PIN Mout_addr_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.984 0.084 22.008 ;
    END
  END Mout_addr_ram[14]
  PIN Mout_addr_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 21.024 59.121 21.048 ;
    END
  END Mout_addr_ram[15]
  PIN Mout_addr_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24.096 59.121 24.12 ;
    END
  END Mout_addr_ram[16]
  PIN Mout_addr_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 21.408 59.121 21.432 ;
    END
  END Mout_addr_ram[17]
  PIN Mout_addr_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 21.504 59.121 21.528 ;
    END
  END Mout_addr_ram[18]
  PIN Mout_addr_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 20.928 59.121 20.952 ;
    END
  END Mout_addr_ram[19]
  PIN Mout_addr_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 27.168 59.121 27.192 ;
    END
  END Mout_addr_ram[1]
  PIN Mout_addr_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 21.792 59.121 21.816 ;
    END
  END Mout_addr_ram[20]
  PIN Mout_addr_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.712 59.121 23.736 ;
    END
  END Mout_addr_ram[21]
  PIN Mout_addr_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 22.656 59.121 22.68 ;
    END
  END Mout_addr_ram[22]
  PIN Mout_addr_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.624 59.037 30.648 59.121 ;
    END
  END Mout_addr_ram[23]
  PIN Mout_addr_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.432 59.037 30.456 59.121 ;
    END
  END Mout_addr_ram[24]
  PIN Mout_addr_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.144 59.037 30.168 59.121 ;
    END
  END Mout_addr_ram[25]
  PIN Mout_addr_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.872 59.037 31.896 59.121 ;
    END
  END Mout_addr_ram[26]
  PIN Mout_addr_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.72 59.037 30.744 59.121 ;
    END
  END Mout_addr_ram[27]
  PIN Mout_addr_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.392 59.037 31.416 59.121 ;
    END
  END Mout_addr_ram[28]
  PIN Mout_addr_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.816 59.037 30.84 59.121 ;
    END
  END Mout_addr_ram[29]
  PIN Mout_addr_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.232 0.084 23.256 ;
    END
  END Mout_addr_ram[2]
  PIN Mout_addr_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.048 59.037 30.072 59.121 ;
    END
  END Mout_addr_ram[30]
  PIN Mout_addr_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.952 59.037 29.976 59.121 ;
    END
  END Mout_addr_ram[31]
  PIN Mout_addr_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.584 59.037 31.608 59.121 ;
    END
  END Mout_addr_ram[32]
  PIN Mout_addr_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.488 59.037 31.512 59.121 ;
    END
  END Mout_addr_ram[33]
  PIN Mout_addr_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.68 59.037 31.704 59.121 ;
    END
  END Mout_addr_ram[34]
  PIN Mout_addr_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.736 59.037 32.76 59.121 ;
    END
  END Mout_addr_ram[35]
  PIN Mout_addr_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.256 59.037 32.28 59.121 ;
    END
  END Mout_addr_ram[36]
  PIN Mout_addr_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.64 59.037 32.664 59.121 ;
    END
  END Mout_addr_ram[37]
  PIN Mout_addr_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.056 59.037 37.08 59.121 ;
    END
  END Mout_addr_ram[38]
  PIN Mout_addr_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.096 59.037 36.12 59.121 ;
    END
  END Mout_addr_ram[39]
  PIN Mout_addr_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.04 0.084 23.064 ;
    END
  END Mout_addr_ram[3]
  PIN Mout_addr_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.424 59.037 35.448 59.121 ;
    END
  END Mout_addr_ram[40]
  PIN Mout_addr_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36 59.037 36.024 59.121 ;
    END
  END Mout_addr_ram[41]
  PIN Mout_addr_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.152 59.037 37.176 59.121 ;
    END
  END Mout_addr_ram[42]
  PIN Mout_addr_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.248 59.037 37.272 59.121 ;
    END
  END Mout_addr_ram[43]
  PIN Mout_addr_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.344 59.037 37.368 59.121 ;
    END
  END Mout_addr_ram[44]
  PIN Mout_addr_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  37.44 59.037 37.464 59.121 ;
    END
  END Mout_addr_ram[45]
  PIN Mout_addr_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.728 0.084 25.752 ;
    END
  END Mout_addr_ram[4]
  PIN Mout_addr_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.248 0.084 25.272 ;
    END
  END Mout_addr_ram[5]
  PIN Mout_addr_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.576 0.084 24.6 ;
    END
  END Mout_addr_ram[6]
  PIN Mout_addr_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.768 0.084 24.792 ;
    END
  END Mout_addr_ram[7]
  PIN Mout_addr_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24 0.084 24.024 ;
    END
  END Mout_addr_ram[8]
  PIN Mout_addr_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.712 0.084 23.736 ;
    END
  END Mout_addr_ram[9]
  PIN Mout_data_ram_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.08 0.084 22.104 ;
    END
  END Mout_data_ram_size[0]
  PIN Mout_data_ram_size[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.568 59.037 29.592 59.121 ;
    END
  END Mout_data_ram_size[10]
  PIN Mout_data_ram_size[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.992 59.037 29.016 59.121 ;
    END
  END Mout_data_ram_size[11]
  PIN Mout_data_ram_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.464 0.084 22.488 ;
    END
  END Mout_data_ram_size[1]
  PIN Mout_data_ram_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.176 0.084 22.2 ;
    END
  END Mout_data_ram_size[2]
  PIN Mout_data_ram_size[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.272 0.084 22.296 ;
    END
  END Mout_data_ram_size[3]
  PIN Mout_data_ram_size[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.656 0.084 22.68 ;
    END
  END Mout_data_ram_size[4]
  PIN Mout_data_ram_size[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24.192 59.121 24.216 ;
    END
  END Mout_data_ram_size[5]
  PIN Mout_data_ram_size[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.472 59.037 29.496 59.121 ;
    END
  END Mout_data_ram_size[6]
  PIN Mout_data_ram_size[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.664 59.037 29.688 59.121 ;
    END
  END Mout_data_ram_size[7]
  PIN Mout_data_ram_size[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.376 59.037 29.4 59.121 ;
    END
  END Mout_data_ram_size[8]
  PIN Mout_data_ram_size[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.76 59.037 29.784 59.121 ;
    END
  END Mout_data_ram_size[9]
  PIN Mout_oe_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.328 59.121 23.352 ;
    END
  END Mout_oe_ram[0]
  PIN Mout_oe_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  35.712 59.037 35.736 59.121 ;
    END
  END Mout_oe_ram[1]
  PIN Mout_we_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 27.84 59.121 27.864 ;
    END
  END Mout_we_ram[0]
  PIN Mout_we_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.28 59.037 29.304 59.121 ;
    END
  END Mout_we_ram[1]
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  54.912 59.037 54.936 59.121 ;
    END
  END clock
  PIN done_port
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.784 0.084 14.808 ;
    END
  END done_port
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.224 59.037 28.248 59.121 ;
    END
  END reset
  PIN start_port
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.168 0 39.192 0.084 ;
    END
  END start_port
  PIN vargs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 26.496 59.121 26.52 ;
    END
  END vargs[0]
  PIN vargs[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 22.56 59.121 22.584 ;
    END
  END vargs[10]
  PIN vargs[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.904 59.121 23.928 ;
    END
  END vargs[11]
  PIN vargs[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 22.944 59.121 22.968 ;
    END
  END vargs[12]
  PIN vargs[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.552 0 39.576 0.084 ;
    END
  END vargs[13]
  PIN vargs[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.84 0 39.864 0.084 ;
    END
  END vargs[14]
  PIN vargs[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.36 0 39.384 0.084 ;
    END
  END vargs[15]
  PIN vargs[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.072 0 39.096 0.084 ;
    END
  END vargs[16]
  PIN vargs[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.472 0 41.496 0.084 ;
    END
  END vargs[17]
  PIN vargs[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.456 0 39.48 0.084 ;
    END
  END vargs[18]
  PIN vargs[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.992 0 41.016 0.084 ;
    END
  END vargs[19]
  PIN vargs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 26.592 59.121 26.616 ;
    END
  END vargs[1]
  PIN vargs[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.8 0 40.824 0.084 ;
    END
  END vargs[20]
  PIN vargs[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.704 0 40.728 0.084 ;
    END
  END vargs[21]
  PIN vargs[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  41.856 0 41.88 0.084 ;
    END
  END vargs[22]
  PIN vargs[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  48.192 0 48.216 0.084 ;
    END
  END vargs[23]
  PIN vargs[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  48.672 0 48.696 0.084 ;
    END
  END vargs[24]
  PIN vargs[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 19.872 59.121 19.896 ;
    END
  END vargs[25]
  PIN vargs[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 21.888 59.121 21.912 ;
    END
  END vargs[26]
  PIN vargs[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.424 59.121 23.448 ;
    END
  END vargs[27]
  PIN vargs[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.52 59.121 23.544 ;
    END
  END vargs[28]
  PIN vargs[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24 59.121 24.024 ;
    END
  END vargs[29]
  PIN vargs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 26.016 59.121 26.04 ;
    END
  END vargs[2]
  PIN vargs[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.808 59.121 23.832 ;
    END
  END vargs[30]
  PIN vargs[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 25.536 59.121 25.56 ;
    END
  END vargs[31]
  PIN vargs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.264 0 39.288 0.084 ;
    END
  END vargs[3]
  PIN vargs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 25.92 59.121 25.944 ;
    END
  END vargs[4]
  PIN vargs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24.864 59.121 24.888 ;
    END
  END vargs[5]
  PIN vargs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24.288 59.121 24.312 ;
    END
  END vargs[6]
  PIN vargs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.616 59.121 23.64 ;
    END
  END vargs[7]
  PIN vargs[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 24.768 59.121 24.792 ;
    END
  END vargs[8]
  PIN vargs[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  59.037 23.04 59.121 23.064 ;
    END
  END vargs[9]
  OBS
    LAYER M1 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M2 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M3 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M4 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M5 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M6 ;
     RECT  0 0 59.121 59.121 ;
    LAYER M7 ;
     RECT  0 0 59.121 59.121 ;
  END
END run_benchmark
END LIBRARY
