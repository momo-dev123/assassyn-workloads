VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA PE_via1_2_3996_18_1_111_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 111 ;
END PE_via1_2_3996_18_1_111_36_36

VIA PE_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END PE_VIA23_1_3_36_36

VIA PE_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END PE_VIA34_1_2_58_52

VIA PE_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END PE_VIA45_1_2_58_58

MACRO PE
  FOREIGN PE 0 0 ;
  CLASS BLOCK ;
  SIZE 6.04 BY 6.04 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  1.458 1.327 1.578 4.613 ;
      LAYER M2 ;
        RECT  1.026 4.581 5.022 4.599 ;
        RECT  1.026 4.041 5.022 4.059 ;
        RECT  1.026 3.501 5.022 3.519 ;
        RECT  1.026 2.961 5.022 2.979 ;
        RECT  1.026 2.421 5.022 2.439 ;
        RECT  1.026 1.881 5.022 1.899 ;
        RECT  1.026 1.341 5.022 1.359 ;
      LAYER M1 ;
        RECT  1.026 4.581 5.022 4.599 ;
        RECT  1.026 4.041 5.022 4.059 ;
        RECT  1.026 3.501 5.022 3.519 ;
        RECT  1.026 2.961 5.022 2.979 ;
        RECT  1.026 2.421 5.022 2.439 ;
        RECT  1.026 1.881 5.022 1.899 ;
        RECT  1.026 1.341 5.022 1.359 ;
      VIA 1.518 4.59 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 PE_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 PE_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 PE_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 PE_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 PE_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 PE_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 PE_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 PE_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 PE_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 PE_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 PE_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 PE_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 PE_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 PE_VIA23_1_3_36_36 ;
      VIA 3.024 4.59 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 4.05 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 3.51 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 2.97 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 2.43 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 1.89 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 1.35 PE_via1_2_3996_18_1_111_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  1.266 1.057 1.386 4.883 ;
      LAYER M2 ;
        RECT  1.026 4.851 5.022 4.869 ;
        RECT  1.026 4.311 5.022 4.329 ;
        RECT  1.026 3.771 5.022 3.789 ;
        RECT  1.026 3.231 5.022 3.249 ;
        RECT  1.026 2.691 5.022 2.709 ;
        RECT  1.026 2.151 5.022 2.169 ;
        RECT  1.026 1.611 5.022 1.629 ;
        RECT  1.026 1.071 5.022 1.089 ;
      LAYER M1 ;
        RECT  1.026 4.851 5.022 4.869 ;
        RECT  1.026 4.311 5.022 4.329 ;
        RECT  1.026 3.771 5.022 3.789 ;
        RECT  1.026 3.231 5.022 3.249 ;
        RECT  1.026 2.691 5.022 2.709 ;
        RECT  1.026 2.151 5.022 2.169 ;
        RECT  1.026 1.611 5.022 1.629 ;
        RECT  1.026 1.071 5.022 1.089 ;
      VIA 1.326 4.86 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 PE_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 PE_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 PE_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 PE_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 PE_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 PE_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 PE_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 PE_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 PE_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 PE_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 PE_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 PE_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 PE_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 PE_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 PE_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 PE_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 PE_VIA23_1_3_36_36 ;
      VIA 3.024 4.86 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 4.32 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 3.78 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 3.24 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 2.7 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 2.16 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 1.62 PE_via1_2_3996_18_1_111_36_36 ;
      VIA 3.024 1.08 PE_via1_2_3996_18_1_111_36_36 ;
    END
  END VSS
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.84 0.084 3.864 ;
    END
  END clock
  PIN io_dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.168 0.084 3.192 ;
    END
  END io_dir
  PIN io_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.728 0 1.752 0.084 ;
    END
  END io_en
  PIN io_inD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.688 0 2.712 0.084 ;
    END
  END io_inD[0]
  PIN io_inD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.168 5.956 3.192 6.04 ;
    END
  END io_inD[1]
  PIN io_inD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.264 0.084 3.288 ;
    END
  END io_inD[2]
  PIN io_inD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.36 0.084 3.384 ;
    END
  END io_inD[3]
  PIN io_inD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.168 0 3.192 0.084 ;
    END
  END io_inD[4]
  PIN io_inD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.688 0.084 2.712 ;
    END
  END io_inD[5]
  PIN io_inD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.112 0.084 2.136 ;
    END
  END io_inD[6]
  PIN io_inD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.264 0 3.288 0.084 ;
    END
  END io_inD[7]
  PIN io_inR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.592 0 2.616 0.084 ;
    END
  END io_inR[0]
  PIN io_inR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 3.36 6.04 3.384 ;
    END
  END io_inR[1]
  PIN io_inR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.456 0.084 3.48 ;
    END
  END io_inR[2]
  PIN io_inR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.688 5.956 2.712 6.04 ;
    END
  END io_inR[3]
  PIN io_inR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 2.784 6.04 2.808 ;
    END
  END io_inR[4]
  PIN io_inR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.592 0.084 2.616 ;
    END
  END io_inR[5]
  PIN io_inR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.016 0.084 2.04 ;
    END
  END io_inR[6]
  PIN io_inR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.456 0 3.48 0.084 ;
    END
  END io_inR[7]
  PIN io_outL[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.552 0 3.576 0.084 ;
    END
  END io_outL[0]
  PIN io_outL[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 3.552 6.04 3.576 ;
    END
  END io_outL[1]
  PIN io_outL[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.648 0.084 3.672 ;
    END
  END io_outL[2]
  PIN io_outL[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.552 5.956 3.576 6.04 ;
    END
  END io_outL[3]
  PIN io_outL[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 2.688 6.04 2.712 ;
    END
  END io_outL[4]
  PIN io_outL[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.784 0 2.808 0.084 ;
    END
  END io_outL[5]
  PIN io_outL[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.304 0 2.328 0.084 ;
    END
  END io_outL[6]
  PIN io_outL[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 2.016 6.04 2.04 ;
    END
  END io_outL[7]
  PIN io_outU[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.744 0 3.768 0.084 ;
    END
  END io_outU[0]
  PIN io_outU[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 3.648 6.04 3.672 ;
    END
  END io_outU[1]
  PIN io_outU[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.744 0.084 3.768 ;
    END
  END io_outU[2]
  PIN io_outU[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.744 5.956 3.768 6.04 ;
    END
  END io_outU[3]
  PIN io_outU[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 2.88 6.04 2.904 ;
    END
  END io_outU[4]
  PIN io_outU[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.976 0 3 0.084 ;
    END
  END io_outU[5]
  PIN io_outU[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.496 0 2.52 0.084 ;
    END
  END io_outU[6]
  PIN io_outU[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.956 2.112 6.04 2.136 ;
    END
  END io_outU[7]
  OBS
    LAYER M1 ;
     RECT  0 0 6.04 6.04 ;
    LAYER M2 ;
     RECT  0 0 6.04 6.04 ;
    LAYER M3 ;
     RECT  0 0 6.04 6.04 ;
    LAYER M4 ;
     RECT  0 0 6.04 6.04 ;
    LAYER M5 ;
     RECT  0 0 6.04 6.04 ;
  END
END PE
END LIBRARY
