VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA run_benchmark_via1_2_39258_18_1_1090_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 1090 ;
END run_benchmark_via1_2_39258_18_1_1090_36_36

VIA run_benchmark_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END run_benchmark_VIA23_1_3_36_36

VIA run_benchmark_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END run_benchmark_VIA34_1_2_58_52

VIA run_benchmark_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END run_benchmark_VIA45_1_2_58_58

VIA run_benchmark_via5_6_120_288_1_2_58_322
  VIARULE M6_M5widePWR1p152 ;
  CUTSIZE 0.024 0.288 ;
  LAYERS M5 V5 M6 ;
  CUTSPACING 0.034 0.034 ;
  ENCLOSURE 0.019 0 0 0 ;
  ROWCOL 1 2 ;
END run_benchmark_via5_6_120_288_1_2_58_322

MACRO run_benchmark
  FOREIGN run_benchmark 0 0 ;
  CLASS BLOCK ;
  SIZE 41.319 BY 41.319 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.458 37.833 37.002 38.121 ;
        RECT  1.458 31.833 37.002 32.121 ;
        RECT  1.458 25.833 37.002 26.121 ;
        RECT  1.458 19.833 37.002 20.121 ;
        RECT  1.458 13.833 37.002 14.121 ;
        RECT  1.458 7.833 37.002 8.121 ;
        RECT  1.458 1.833 37.002 2.121 ;
      LAYER M5 ;
        RECT  36.882 1.327 37.002 40.253 ;
        RECT  30.978 1.327 31.098 40.253 ;
        RECT  25.074 1.327 25.194 40.253 ;
        RECT  19.17 1.327 19.29 40.253 ;
        RECT  13.266 1.327 13.386 40.253 ;
        RECT  7.362 1.327 7.482 40.253 ;
        RECT  1.458 1.327 1.578 40.253 ;
      LAYER M2 ;
        RECT  1.026 40.221 40.284 40.239 ;
        RECT  1.026 39.681 40.284 39.699 ;
        RECT  1.026 39.141 40.284 39.159 ;
        RECT  1.026 38.601 40.284 38.619 ;
        RECT  1.026 38.061 40.284 38.079 ;
        RECT  1.026 37.521 40.284 37.539 ;
        RECT  1.026 36.981 40.284 36.999 ;
        RECT  1.026 36.441 40.284 36.459 ;
        RECT  1.026 35.901 40.284 35.919 ;
        RECT  1.026 35.361 40.284 35.379 ;
        RECT  1.026 34.821 40.284 34.839 ;
        RECT  1.026 34.281 40.284 34.299 ;
        RECT  1.026 33.741 40.284 33.759 ;
        RECT  1.026 33.201 40.284 33.219 ;
        RECT  1.026 32.661 40.284 32.679 ;
        RECT  1.026 32.121 40.284 32.139 ;
        RECT  1.026 31.581 40.284 31.599 ;
        RECT  1.026 31.041 40.284 31.059 ;
        RECT  1.026 30.501 40.284 30.519 ;
        RECT  1.026 29.961 40.284 29.979 ;
        RECT  1.026 29.421 40.284 29.439 ;
        RECT  1.026 28.881 40.284 28.899 ;
        RECT  1.026 28.341 40.284 28.359 ;
        RECT  1.026 27.801 40.284 27.819 ;
        RECT  1.026 27.261 40.284 27.279 ;
        RECT  1.026 26.721 40.284 26.739 ;
        RECT  1.026 26.181 40.284 26.199 ;
        RECT  1.026 25.641 40.284 25.659 ;
        RECT  1.026 25.101 40.284 25.119 ;
        RECT  1.026 24.561 40.284 24.579 ;
        RECT  1.026 24.021 40.284 24.039 ;
        RECT  1.026 23.481 40.284 23.499 ;
        RECT  1.026 22.941 40.284 22.959 ;
        RECT  1.026 22.401 40.284 22.419 ;
        RECT  1.026 21.861 40.284 21.879 ;
        RECT  1.026 21.321 40.284 21.339 ;
        RECT  1.026 20.781 40.284 20.799 ;
        RECT  1.026 20.241 40.284 20.259 ;
        RECT  1.026 19.701 40.284 19.719 ;
        RECT  1.026 19.161 40.284 19.179 ;
        RECT  1.026 18.621 40.284 18.639 ;
        RECT  1.026 18.081 40.284 18.099 ;
        RECT  1.026 17.541 40.284 17.559 ;
        RECT  1.026 17.001 40.284 17.019 ;
        RECT  1.026 16.461 40.284 16.479 ;
        RECT  1.026 15.921 40.284 15.939 ;
        RECT  1.026 15.381 40.284 15.399 ;
        RECT  1.026 14.841 40.284 14.859 ;
        RECT  1.026 14.301 40.284 14.319 ;
        RECT  1.026 13.761 40.284 13.779 ;
        RECT  1.026 13.221 40.284 13.239 ;
        RECT  1.026 12.681 40.284 12.699 ;
        RECT  1.026 12.141 40.284 12.159 ;
        RECT  1.026 11.601 40.284 11.619 ;
        RECT  1.026 11.061 40.284 11.079 ;
        RECT  1.026 10.521 40.284 10.539 ;
        RECT  1.026 9.981 40.284 9.999 ;
        RECT  1.026 9.441 40.284 9.459 ;
        RECT  1.026 8.901 40.284 8.919 ;
        RECT  1.026 8.361 40.284 8.379 ;
        RECT  1.026 7.821 40.284 7.839 ;
        RECT  1.026 7.281 40.284 7.299 ;
        RECT  1.026 6.741 40.284 6.759 ;
        RECT  1.026 6.201 40.284 6.219 ;
        RECT  1.026 5.661 40.284 5.679 ;
        RECT  1.026 5.121 40.284 5.139 ;
        RECT  1.026 4.581 40.284 4.599 ;
        RECT  1.026 4.041 40.284 4.059 ;
        RECT  1.026 3.501 40.284 3.519 ;
        RECT  1.026 2.961 40.284 2.979 ;
        RECT  1.026 2.421 40.284 2.439 ;
        RECT  1.026 1.881 40.284 1.899 ;
        RECT  1.026 1.341 40.284 1.359 ;
      LAYER M1 ;
        RECT  1.026 40.221 40.284 40.239 ;
        RECT  1.026 39.681 40.284 39.699 ;
        RECT  1.026 39.141 40.284 39.159 ;
        RECT  1.026 38.601 40.284 38.619 ;
        RECT  1.026 38.061 40.284 38.079 ;
        RECT  1.026 37.521 40.284 37.539 ;
        RECT  1.026 36.981 40.284 36.999 ;
        RECT  1.026 36.441 40.284 36.459 ;
        RECT  1.026 35.901 40.284 35.919 ;
        RECT  1.026 35.361 40.284 35.379 ;
        RECT  1.026 34.821 40.284 34.839 ;
        RECT  1.026 34.281 40.284 34.299 ;
        RECT  1.026 33.741 40.284 33.759 ;
        RECT  1.026 33.201 40.284 33.219 ;
        RECT  1.026 32.661 40.284 32.679 ;
        RECT  1.026 32.121 40.284 32.139 ;
        RECT  1.026 31.581 40.284 31.599 ;
        RECT  1.026 31.041 40.284 31.059 ;
        RECT  1.026 30.501 40.284 30.519 ;
        RECT  1.026 29.961 40.284 29.979 ;
        RECT  1.026 29.421 40.284 29.439 ;
        RECT  1.026 28.881 40.284 28.899 ;
        RECT  1.026 28.341 40.284 28.359 ;
        RECT  1.026 27.801 40.284 27.819 ;
        RECT  1.026 27.261 40.284 27.279 ;
        RECT  1.026 26.721 40.284 26.739 ;
        RECT  1.026 26.181 40.284 26.199 ;
        RECT  1.026 25.641 40.284 25.659 ;
        RECT  1.026 25.101 40.284 25.119 ;
        RECT  1.026 24.561 40.284 24.579 ;
        RECT  1.026 24.021 40.284 24.039 ;
        RECT  1.026 23.481 40.284 23.499 ;
        RECT  1.026 22.941 40.284 22.959 ;
        RECT  1.026 22.401 40.284 22.419 ;
        RECT  1.026 21.861 40.284 21.879 ;
        RECT  1.026 21.321 40.284 21.339 ;
        RECT  1.026 20.781 40.284 20.799 ;
        RECT  1.026 20.241 40.284 20.259 ;
        RECT  1.026 19.701 40.284 19.719 ;
        RECT  1.026 19.161 40.284 19.179 ;
        RECT  1.026 18.621 40.284 18.639 ;
        RECT  1.026 18.081 40.284 18.099 ;
        RECT  1.026 17.541 40.284 17.559 ;
        RECT  1.026 17.001 40.284 17.019 ;
        RECT  1.026 16.461 40.284 16.479 ;
        RECT  1.026 15.921 40.284 15.939 ;
        RECT  1.026 15.381 40.284 15.399 ;
        RECT  1.026 14.841 40.284 14.859 ;
        RECT  1.026 14.301 40.284 14.319 ;
        RECT  1.026 13.761 40.284 13.779 ;
        RECT  1.026 13.221 40.284 13.239 ;
        RECT  1.026 12.681 40.284 12.699 ;
        RECT  1.026 12.141 40.284 12.159 ;
        RECT  1.026 11.601 40.284 11.619 ;
        RECT  1.026 11.061 40.284 11.079 ;
        RECT  1.026 10.521 40.284 10.539 ;
        RECT  1.026 9.981 40.284 9.999 ;
        RECT  1.026 9.441 40.284 9.459 ;
        RECT  1.026 8.901 40.284 8.919 ;
        RECT  1.026 8.361 40.284 8.379 ;
        RECT  1.026 7.821 40.284 7.839 ;
        RECT  1.026 7.281 40.284 7.299 ;
        RECT  1.026 6.741 40.284 6.759 ;
        RECT  1.026 6.201 40.284 6.219 ;
        RECT  1.026 5.661 40.284 5.679 ;
        RECT  1.026 5.121 40.284 5.139 ;
        RECT  1.026 4.581 40.284 4.599 ;
        RECT  1.026 4.041 40.284 4.059 ;
        RECT  1.026 3.501 40.284 3.519 ;
        RECT  1.026 2.961 40.284 2.979 ;
        RECT  1.026 2.421 40.284 2.439 ;
        RECT  1.026 1.881 40.284 1.899 ;
        RECT  1.026 1.341 40.284 1.359 ;
      VIA 36.942 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 31.038 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 25.134 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.23 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.326 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 37.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 31.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 25.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 19.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 13.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 7.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 1.977 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.942 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 40.213 36.987 40.247 ;
      VIA 36.942 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.673 36.987 39.707 ;
      VIA 36.942 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 39.133 36.987 39.167 ;
      VIA 36.942 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.593 36.987 38.627 ;
      VIA 36.942 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 38.053 36.987 38.087 ;
      VIA 36.942 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 37.513 36.987 37.547 ;
      VIA 36.942 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.973 36.987 37.007 ;
      VIA 36.942 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 36.433 36.987 36.467 ;
      VIA 36.942 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.893 36.987 35.927 ;
      VIA 36.942 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 35.353 36.987 35.387 ;
      VIA 36.942 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.813 36.987 34.847 ;
      VIA 36.942 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 34.273 36.987 34.307 ;
      VIA 36.942 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.733 36.987 33.767 ;
      VIA 36.942 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 33.193 36.987 33.227 ;
      VIA 36.942 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.653 36.987 32.687 ;
      VIA 36.942 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 32.113 36.987 32.147 ;
      VIA 36.942 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.573 36.987 31.607 ;
      VIA 36.942 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 31.033 36.987 31.067 ;
      VIA 36.942 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 30.493 36.987 30.527 ;
      VIA 36.942 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.953 36.987 29.987 ;
      VIA 36.942 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 29.413 36.987 29.447 ;
      VIA 36.942 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.873 36.987 28.907 ;
      VIA 36.942 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 28.333 36.987 28.367 ;
      VIA 36.942 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.793 36.987 27.827 ;
      VIA 36.942 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 27.253 36.987 27.287 ;
      VIA 36.942 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.713 36.987 26.747 ;
      VIA 36.942 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 26.173 36.987 26.207 ;
      VIA 36.942 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.633 36.987 25.667 ;
      VIA 36.942 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 25.093 36.987 25.127 ;
      VIA 36.942 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.553 36.987 24.587 ;
      VIA 36.942 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 24.013 36.987 24.047 ;
      VIA 36.942 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 23.473 36.987 23.507 ;
      VIA 36.942 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.933 36.987 22.967 ;
      VIA 36.942 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 22.393 36.987 22.427 ;
      VIA 36.942 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.853 36.987 21.887 ;
      VIA 36.942 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 21.313 36.987 21.347 ;
      VIA 36.942 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.773 36.987 20.807 ;
      VIA 36.942 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 20.233 36.987 20.267 ;
      VIA 36.942 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.693 36.987 19.727 ;
      VIA 36.942 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 19.153 36.987 19.187 ;
      VIA 36.942 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.613 36.987 18.647 ;
      VIA 36.942 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 18.073 36.987 18.107 ;
      VIA 36.942 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 17.533 36.987 17.567 ;
      VIA 36.942 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.993 36.987 17.027 ;
      VIA 36.942 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 16.453 36.987 16.487 ;
      VIA 36.942 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.913 36.987 15.947 ;
      VIA 36.942 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 15.373 36.987 15.407 ;
      VIA 36.942 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.833 36.987 14.867 ;
      VIA 36.942 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 14.293 36.987 14.327 ;
      VIA 36.942 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.753 36.987 13.787 ;
      VIA 36.942 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 13.213 36.987 13.247 ;
      VIA 36.942 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.673 36.987 12.707 ;
      VIA 36.942 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 12.133 36.987 12.167 ;
      VIA 36.942 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.593 36.987 11.627 ;
      VIA 36.942 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 11.053 36.987 11.087 ;
      VIA 36.942 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 10.513 36.987 10.547 ;
      VIA 36.942 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.973 36.987 10.007 ;
      VIA 36.942 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 9.433 36.987 9.467 ;
      VIA 36.942 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.893 36.987 8.927 ;
      VIA 36.942 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 8.353 36.987 8.387 ;
      VIA 36.942 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.813 36.987 7.847 ;
      VIA 36.942 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 7.273 36.987 7.307 ;
      VIA 36.942 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.733 36.987 6.767 ;
      VIA 36.942 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 6.193 36.987 6.227 ;
      VIA 36.942 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.653 36.987 5.687 ;
      VIA 36.942 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 5.113 36.987 5.147 ;
      VIA 36.942 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.573 36.987 4.607 ;
      VIA 36.942 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 4.033 36.987 4.067 ;
      VIA 36.942 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 3.493 36.987 3.527 ;
      VIA 36.942 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.953 36.987 2.987 ;
      VIA 36.942 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 2.413 36.987 2.447 ;
      VIA 36.942 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.873 36.987 1.907 ;
      VIA 36.942 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.942 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.897 1.333 36.987 1.367 ;
      VIA 36.942 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.942 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 40.213 31.083 40.247 ;
      VIA 31.038 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.673 31.083 39.707 ;
      VIA 31.038 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 39.133 31.083 39.167 ;
      VIA 31.038 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.593 31.083 38.627 ;
      VIA 31.038 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 38.053 31.083 38.087 ;
      VIA 31.038 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 37.513 31.083 37.547 ;
      VIA 31.038 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.973 31.083 37.007 ;
      VIA 31.038 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 36.433 31.083 36.467 ;
      VIA 31.038 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.893 31.083 35.927 ;
      VIA 31.038 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 35.353 31.083 35.387 ;
      VIA 31.038 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.813 31.083 34.847 ;
      VIA 31.038 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 34.273 31.083 34.307 ;
      VIA 31.038 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.733 31.083 33.767 ;
      VIA 31.038 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 33.193 31.083 33.227 ;
      VIA 31.038 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.653 31.083 32.687 ;
      VIA 31.038 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 32.113 31.083 32.147 ;
      VIA 31.038 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.573 31.083 31.607 ;
      VIA 31.038 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 31.033 31.083 31.067 ;
      VIA 31.038 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 30.493 31.083 30.527 ;
      VIA 31.038 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.953 31.083 29.987 ;
      VIA 31.038 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 29.413 31.083 29.447 ;
      VIA 31.038 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.873 31.083 28.907 ;
      VIA 31.038 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 28.333 31.083 28.367 ;
      VIA 31.038 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.793 31.083 27.827 ;
      VIA 31.038 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 27.253 31.083 27.287 ;
      VIA 31.038 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.713 31.083 26.747 ;
      VIA 31.038 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 26.173 31.083 26.207 ;
      VIA 31.038 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.633 31.083 25.667 ;
      VIA 31.038 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 25.093 31.083 25.127 ;
      VIA 31.038 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.553 31.083 24.587 ;
      VIA 31.038 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 24.013 31.083 24.047 ;
      VIA 31.038 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 23.473 31.083 23.507 ;
      VIA 31.038 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.933 31.083 22.967 ;
      VIA 31.038 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 22.393 31.083 22.427 ;
      VIA 31.038 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.853 31.083 21.887 ;
      VIA 31.038 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 21.313 31.083 21.347 ;
      VIA 31.038 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.773 31.083 20.807 ;
      VIA 31.038 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 20.233 31.083 20.267 ;
      VIA 31.038 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.693 31.083 19.727 ;
      VIA 31.038 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 19.153 31.083 19.187 ;
      VIA 31.038 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.613 31.083 18.647 ;
      VIA 31.038 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 18.073 31.083 18.107 ;
      VIA 31.038 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 17.533 31.083 17.567 ;
      VIA 31.038 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.993 31.083 17.027 ;
      VIA 31.038 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 16.453 31.083 16.487 ;
      VIA 31.038 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.913 31.083 15.947 ;
      VIA 31.038 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 15.373 31.083 15.407 ;
      VIA 31.038 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.833 31.083 14.867 ;
      VIA 31.038 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 14.293 31.083 14.327 ;
      VIA 31.038 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.753 31.083 13.787 ;
      VIA 31.038 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 13.213 31.083 13.247 ;
      VIA 31.038 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.673 31.083 12.707 ;
      VIA 31.038 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 12.133 31.083 12.167 ;
      VIA 31.038 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.593 31.083 11.627 ;
      VIA 31.038 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 11.053 31.083 11.087 ;
      VIA 31.038 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 10.513 31.083 10.547 ;
      VIA 31.038 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.973 31.083 10.007 ;
      VIA 31.038 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 9.433 31.083 9.467 ;
      VIA 31.038 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.893 31.083 8.927 ;
      VIA 31.038 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 8.353 31.083 8.387 ;
      VIA 31.038 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.813 31.083 7.847 ;
      VIA 31.038 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 7.273 31.083 7.307 ;
      VIA 31.038 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.733 31.083 6.767 ;
      VIA 31.038 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 6.193 31.083 6.227 ;
      VIA 31.038 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.653 31.083 5.687 ;
      VIA 31.038 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 5.113 31.083 5.147 ;
      VIA 31.038 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.573 31.083 4.607 ;
      VIA 31.038 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 4.033 31.083 4.067 ;
      VIA 31.038 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 3.493 31.083 3.527 ;
      VIA 31.038 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.953 31.083 2.987 ;
      VIA 31.038 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 2.413 31.083 2.447 ;
      VIA 31.038 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.873 31.083 1.907 ;
      VIA 31.038 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 31.038 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.993 1.333 31.083 1.367 ;
      VIA 31.038 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 31.038 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 40.213 25.179 40.247 ;
      VIA 25.134 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.673 25.179 39.707 ;
      VIA 25.134 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 39.133 25.179 39.167 ;
      VIA 25.134 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.593 25.179 38.627 ;
      VIA 25.134 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 38.053 25.179 38.087 ;
      VIA 25.134 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 37.513 25.179 37.547 ;
      VIA 25.134 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.973 25.179 37.007 ;
      VIA 25.134 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 36.433 25.179 36.467 ;
      VIA 25.134 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.893 25.179 35.927 ;
      VIA 25.134 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 35.353 25.179 35.387 ;
      VIA 25.134 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.813 25.179 34.847 ;
      VIA 25.134 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 34.273 25.179 34.307 ;
      VIA 25.134 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.733 25.179 33.767 ;
      VIA 25.134 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 33.193 25.179 33.227 ;
      VIA 25.134 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.653 25.179 32.687 ;
      VIA 25.134 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 32.113 25.179 32.147 ;
      VIA 25.134 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.573 25.179 31.607 ;
      VIA 25.134 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 31.033 25.179 31.067 ;
      VIA 25.134 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 30.493 25.179 30.527 ;
      VIA 25.134 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.953 25.179 29.987 ;
      VIA 25.134 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 29.413 25.179 29.447 ;
      VIA 25.134 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.873 25.179 28.907 ;
      VIA 25.134 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 28.333 25.179 28.367 ;
      VIA 25.134 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.793 25.179 27.827 ;
      VIA 25.134 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 27.253 25.179 27.287 ;
      VIA 25.134 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.713 25.179 26.747 ;
      VIA 25.134 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 26.173 25.179 26.207 ;
      VIA 25.134 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.633 25.179 25.667 ;
      VIA 25.134 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 25.093 25.179 25.127 ;
      VIA 25.134 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.553 25.179 24.587 ;
      VIA 25.134 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 24.013 25.179 24.047 ;
      VIA 25.134 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 23.473 25.179 23.507 ;
      VIA 25.134 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.933 25.179 22.967 ;
      VIA 25.134 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 22.393 25.179 22.427 ;
      VIA 25.134 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.853 25.179 21.887 ;
      VIA 25.134 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 21.313 25.179 21.347 ;
      VIA 25.134 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.773 25.179 20.807 ;
      VIA 25.134 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 20.233 25.179 20.267 ;
      VIA 25.134 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.693 25.179 19.727 ;
      VIA 25.134 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 19.153 25.179 19.187 ;
      VIA 25.134 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.613 25.179 18.647 ;
      VIA 25.134 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 18.073 25.179 18.107 ;
      VIA 25.134 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 17.533 25.179 17.567 ;
      VIA 25.134 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.993 25.179 17.027 ;
      VIA 25.134 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 16.453 25.179 16.487 ;
      VIA 25.134 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.913 25.179 15.947 ;
      VIA 25.134 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 15.373 25.179 15.407 ;
      VIA 25.134 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.833 25.179 14.867 ;
      VIA 25.134 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 14.293 25.179 14.327 ;
      VIA 25.134 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.753 25.179 13.787 ;
      VIA 25.134 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 13.213 25.179 13.247 ;
      VIA 25.134 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.673 25.179 12.707 ;
      VIA 25.134 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 12.133 25.179 12.167 ;
      VIA 25.134 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.593 25.179 11.627 ;
      VIA 25.134 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 11.053 25.179 11.087 ;
      VIA 25.134 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 10.513 25.179 10.547 ;
      VIA 25.134 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.973 25.179 10.007 ;
      VIA 25.134 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 9.433 25.179 9.467 ;
      VIA 25.134 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.893 25.179 8.927 ;
      VIA 25.134 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 8.353 25.179 8.387 ;
      VIA 25.134 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.813 25.179 7.847 ;
      VIA 25.134 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 7.273 25.179 7.307 ;
      VIA 25.134 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.733 25.179 6.767 ;
      VIA 25.134 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 6.193 25.179 6.227 ;
      VIA 25.134 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.653 25.179 5.687 ;
      VIA 25.134 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 5.113 25.179 5.147 ;
      VIA 25.134 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.573 25.179 4.607 ;
      VIA 25.134 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 4.033 25.179 4.067 ;
      VIA 25.134 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 3.493 25.179 3.527 ;
      VIA 25.134 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.953 25.179 2.987 ;
      VIA 25.134 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 2.413 25.179 2.447 ;
      VIA 25.134 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.873 25.179 1.907 ;
      VIA 25.134 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 25.134 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  25.089 1.333 25.179 1.367 ;
      VIA 25.134 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 25.134 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 40.213 19.275 40.247 ;
      VIA 19.23 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.673 19.275 39.707 ;
      VIA 19.23 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 39.133 19.275 39.167 ;
      VIA 19.23 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.593 19.275 38.627 ;
      VIA 19.23 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 38.053 19.275 38.087 ;
      VIA 19.23 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 37.513 19.275 37.547 ;
      VIA 19.23 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.973 19.275 37.007 ;
      VIA 19.23 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 36.433 19.275 36.467 ;
      VIA 19.23 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.893 19.275 35.927 ;
      VIA 19.23 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 35.353 19.275 35.387 ;
      VIA 19.23 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.813 19.275 34.847 ;
      VIA 19.23 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 34.273 19.275 34.307 ;
      VIA 19.23 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.733 19.275 33.767 ;
      VIA 19.23 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 33.193 19.275 33.227 ;
      VIA 19.23 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.653 19.275 32.687 ;
      VIA 19.23 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 32.113 19.275 32.147 ;
      VIA 19.23 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.573 19.275 31.607 ;
      VIA 19.23 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 31.033 19.275 31.067 ;
      VIA 19.23 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 30.493 19.275 30.527 ;
      VIA 19.23 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.953 19.275 29.987 ;
      VIA 19.23 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 29.413 19.275 29.447 ;
      VIA 19.23 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.873 19.275 28.907 ;
      VIA 19.23 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 28.333 19.275 28.367 ;
      VIA 19.23 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.793 19.275 27.827 ;
      VIA 19.23 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 27.253 19.275 27.287 ;
      VIA 19.23 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.713 19.275 26.747 ;
      VIA 19.23 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 26.173 19.275 26.207 ;
      VIA 19.23 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.633 19.275 25.667 ;
      VIA 19.23 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 25.093 19.275 25.127 ;
      VIA 19.23 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.553 19.275 24.587 ;
      VIA 19.23 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 24.013 19.275 24.047 ;
      VIA 19.23 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 23.473 19.275 23.507 ;
      VIA 19.23 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.933 19.275 22.967 ;
      VIA 19.23 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 22.393 19.275 22.427 ;
      VIA 19.23 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.853 19.275 21.887 ;
      VIA 19.23 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 21.313 19.275 21.347 ;
      VIA 19.23 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.773 19.275 20.807 ;
      VIA 19.23 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 20.233 19.275 20.267 ;
      VIA 19.23 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.693 19.275 19.727 ;
      VIA 19.23 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 19.153 19.275 19.187 ;
      VIA 19.23 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.613 19.275 18.647 ;
      VIA 19.23 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 18.073 19.275 18.107 ;
      VIA 19.23 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 17.533 19.275 17.567 ;
      VIA 19.23 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.993 19.275 17.027 ;
      VIA 19.23 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 16.453 19.275 16.487 ;
      VIA 19.23 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.913 19.275 15.947 ;
      VIA 19.23 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 15.373 19.275 15.407 ;
      VIA 19.23 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.833 19.275 14.867 ;
      VIA 19.23 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 14.293 19.275 14.327 ;
      VIA 19.23 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.753 19.275 13.787 ;
      VIA 19.23 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 13.213 19.275 13.247 ;
      VIA 19.23 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.673 19.275 12.707 ;
      VIA 19.23 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 12.133 19.275 12.167 ;
      VIA 19.23 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.593 19.275 11.627 ;
      VIA 19.23 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 11.053 19.275 11.087 ;
      VIA 19.23 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 10.513 19.275 10.547 ;
      VIA 19.23 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.973 19.275 10.007 ;
      VIA 19.23 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 9.433 19.275 9.467 ;
      VIA 19.23 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.893 19.275 8.927 ;
      VIA 19.23 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 8.353 19.275 8.387 ;
      VIA 19.23 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.813 19.275 7.847 ;
      VIA 19.23 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 7.273 19.275 7.307 ;
      VIA 19.23 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.733 19.275 6.767 ;
      VIA 19.23 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 6.193 19.275 6.227 ;
      VIA 19.23 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.653 19.275 5.687 ;
      VIA 19.23 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 5.113 19.275 5.147 ;
      VIA 19.23 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.573 19.275 4.607 ;
      VIA 19.23 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 4.033 19.275 4.067 ;
      VIA 19.23 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 3.493 19.275 3.527 ;
      VIA 19.23 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.953 19.275 2.987 ;
      VIA 19.23 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 2.413 19.275 2.447 ;
      VIA 19.23 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.873 19.275 1.907 ;
      VIA 19.23 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.23 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  19.185 1.333 19.275 1.367 ;
      VIA 19.23 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.23 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 40.213 13.371 40.247 ;
      VIA 13.326 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.673 13.371 39.707 ;
      VIA 13.326 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 39.133 13.371 39.167 ;
      VIA 13.326 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.593 13.371 38.627 ;
      VIA 13.326 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 38.053 13.371 38.087 ;
      VIA 13.326 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 37.513 13.371 37.547 ;
      VIA 13.326 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.973 13.371 37.007 ;
      VIA 13.326 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 36.433 13.371 36.467 ;
      VIA 13.326 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.893 13.371 35.927 ;
      VIA 13.326 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 35.353 13.371 35.387 ;
      VIA 13.326 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.813 13.371 34.847 ;
      VIA 13.326 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 34.273 13.371 34.307 ;
      VIA 13.326 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.733 13.371 33.767 ;
      VIA 13.326 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 33.193 13.371 33.227 ;
      VIA 13.326 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.653 13.371 32.687 ;
      VIA 13.326 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 32.113 13.371 32.147 ;
      VIA 13.326 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.573 13.371 31.607 ;
      VIA 13.326 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 31.033 13.371 31.067 ;
      VIA 13.326 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 30.493 13.371 30.527 ;
      VIA 13.326 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.953 13.371 29.987 ;
      VIA 13.326 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 29.413 13.371 29.447 ;
      VIA 13.326 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.873 13.371 28.907 ;
      VIA 13.326 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 28.333 13.371 28.367 ;
      VIA 13.326 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.793 13.371 27.827 ;
      VIA 13.326 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 27.253 13.371 27.287 ;
      VIA 13.326 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.713 13.371 26.747 ;
      VIA 13.326 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 26.173 13.371 26.207 ;
      VIA 13.326 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.633 13.371 25.667 ;
      VIA 13.326 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 25.093 13.371 25.127 ;
      VIA 13.326 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.553 13.371 24.587 ;
      VIA 13.326 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 24.013 13.371 24.047 ;
      VIA 13.326 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 23.473 13.371 23.507 ;
      VIA 13.326 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.933 13.371 22.967 ;
      VIA 13.326 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 22.393 13.371 22.427 ;
      VIA 13.326 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.853 13.371 21.887 ;
      VIA 13.326 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 21.313 13.371 21.347 ;
      VIA 13.326 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.773 13.371 20.807 ;
      VIA 13.326 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 20.233 13.371 20.267 ;
      VIA 13.326 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.693 13.371 19.727 ;
      VIA 13.326 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 19.153 13.371 19.187 ;
      VIA 13.326 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.613 13.371 18.647 ;
      VIA 13.326 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 18.073 13.371 18.107 ;
      VIA 13.326 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 17.533 13.371 17.567 ;
      VIA 13.326 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.993 13.371 17.027 ;
      VIA 13.326 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 16.453 13.371 16.487 ;
      VIA 13.326 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.913 13.371 15.947 ;
      VIA 13.326 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 15.373 13.371 15.407 ;
      VIA 13.326 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.833 13.371 14.867 ;
      VIA 13.326 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 14.293 13.371 14.327 ;
      VIA 13.326 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.753 13.371 13.787 ;
      VIA 13.326 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 13.213 13.371 13.247 ;
      VIA 13.326 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.673 13.371 12.707 ;
      VIA 13.326 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 12.133 13.371 12.167 ;
      VIA 13.326 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.593 13.371 11.627 ;
      VIA 13.326 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 11.053 13.371 11.087 ;
      VIA 13.326 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 10.513 13.371 10.547 ;
      VIA 13.326 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.973 13.371 10.007 ;
      VIA 13.326 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 9.433 13.371 9.467 ;
      VIA 13.326 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.893 13.371 8.927 ;
      VIA 13.326 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 8.353 13.371 8.387 ;
      VIA 13.326 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.813 13.371 7.847 ;
      VIA 13.326 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 7.273 13.371 7.307 ;
      VIA 13.326 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.733 13.371 6.767 ;
      VIA 13.326 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 6.193 13.371 6.227 ;
      VIA 13.326 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.653 13.371 5.687 ;
      VIA 13.326 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 5.113 13.371 5.147 ;
      VIA 13.326 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.573 13.371 4.607 ;
      VIA 13.326 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 4.033 13.371 4.067 ;
      VIA 13.326 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 3.493 13.371 3.527 ;
      VIA 13.326 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.953 13.371 2.987 ;
      VIA 13.326 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 2.413 13.371 2.447 ;
      VIA 13.326 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.873 13.371 1.907 ;
      VIA 13.326 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.326 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.281 1.333 13.371 1.367 ;
      VIA 13.326 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.326 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 40.213 7.467 40.247 ;
      VIA 7.422 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.673 7.467 39.707 ;
      VIA 7.422 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 39.133 7.467 39.167 ;
      VIA 7.422 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.593 7.467 38.627 ;
      VIA 7.422 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 38.053 7.467 38.087 ;
      VIA 7.422 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 37.513 7.467 37.547 ;
      VIA 7.422 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.973 7.467 37.007 ;
      VIA 7.422 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 36.433 7.467 36.467 ;
      VIA 7.422 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.893 7.467 35.927 ;
      VIA 7.422 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 35.353 7.467 35.387 ;
      VIA 7.422 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.813 7.467 34.847 ;
      VIA 7.422 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 34.273 7.467 34.307 ;
      VIA 7.422 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.733 7.467 33.767 ;
      VIA 7.422 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 33.193 7.467 33.227 ;
      VIA 7.422 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.653 7.467 32.687 ;
      VIA 7.422 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 32.113 7.467 32.147 ;
      VIA 7.422 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.573 7.467 31.607 ;
      VIA 7.422 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 31.033 7.467 31.067 ;
      VIA 7.422 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 30.493 7.467 30.527 ;
      VIA 7.422 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.953 7.467 29.987 ;
      VIA 7.422 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 29.413 7.467 29.447 ;
      VIA 7.422 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.873 7.467 28.907 ;
      VIA 7.422 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 28.333 7.467 28.367 ;
      VIA 7.422 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.793 7.467 27.827 ;
      VIA 7.422 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 27.253 7.467 27.287 ;
      VIA 7.422 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.713 7.467 26.747 ;
      VIA 7.422 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 26.173 7.467 26.207 ;
      VIA 7.422 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.633 7.467 25.667 ;
      VIA 7.422 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 25.093 7.467 25.127 ;
      VIA 7.422 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.553 7.467 24.587 ;
      VIA 7.422 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 24.013 7.467 24.047 ;
      VIA 7.422 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 23.473 7.467 23.507 ;
      VIA 7.422 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.933 7.467 22.967 ;
      VIA 7.422 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 22.393 7.467 22.427 ;
      VIA 7.422 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.853 7.467 21.887 ;
      VIA 7.422 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 21.313 7.467 21.347 ;
      VIA 7.422 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.773 7.467 20.807 ;
      VIA 7.422 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 20.233 7.467 20.267 ;
      VIA 7.422 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.693 7.467 19.727 ;
      VIA 7.422 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 19.153 7.467 19.187 ;
      VIA 7.422 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.613 7.467 18.647 ;
      VIA 7.422 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 18.073 7.467 18.107 ;
      VIA 7.422 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 17.533 7.467 17.567 ;
      VIA 7.422 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.993 7.467 17.027 ;
      VIA 7.422 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 16.453 7.467 16.487 ;
      VIA 7.422 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.913 7.467 15.947 ;
      VIA 7.422 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 15.373 7.467 15.407 ;
      VIA 7.422 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.833 7.467 14.867 ;
      VIA 7.422 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 14.293 7.467 14.327 ;
      VIA 7.422 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.753 7.467 13.787 ;
      VIA 7.422 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 13.213 7.467 13.247 ;
      VIA 7.422 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.673 7.467 12.707 ;
      VIA 7.422 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 12.133 7.467 12.167 ;
      VIA 7.422 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.593 7.467 11.627 ;
      VIA 7.422 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.053 7.467 11.087 ;
      VIA 7.422 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 10.513 7.467 10.547 ;
      VIA 7.422 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.973 7.467 10.007 ;
      VIA 7.422 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.433 7.467 9.467 ;
      VIA 7.422 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.893 7.467 8.927 ;
      VIA 7.422 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.353 7.467 8.387 ;
      VIA 7.422 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.813 7.467 7.847 ;
      VIA 7.422 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.273 7.467 7.307 ;
      VIA 7.422 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.733 7.467 6.767 ;
      VIA 7.422 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.193 7.467 6.227 ;
      VIA 7.422 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.653 7.467 5.687 ;
      VIA 7.422 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.113 7.467 5.147 ;
      VIA 7.422 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.573 7.467 4.607 ;
      VIA 7.422 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.033 7.467 4.067 ;
      VIA 7.422 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 3.493 7.467 3.527 ;
      VIA 7.422 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.953 7.467 2.987 ;
      VIA 7.422 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.413 7.467 2.447 ;
      VIA 7.422 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.873 7.467 1.907 ;
      VIA 7.422 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.422 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.333 7.467 1.367 ;
      VIA 7.422 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.422 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 40.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 40.213 1.563 40.247 ;
      VIA 1.518 40.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 40.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.673 1.563 39.707 ;
      VIA 1.518 39.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 39.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 39.133 1.563 39.167 ;
      VIA 1.518 39.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 39.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.593 1.563 38.627 ;
      VIA 1.518 38.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 38.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 38.053 1.563 38.087 ;
      VIA 1.518 38.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 38.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 37.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 37.513 1.563 37.547 ;
      VIA 1.518 37.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 37.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.973 1.563 37.007 ;
      VIA 1.518 36.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 36.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 36.433 1.563 36.467 ;
      VIA 1.518 36.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 36.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.893 1.563 35.927 ;
      VIA 1.518 35.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 35.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 35.353 1.563 35.387 ;
      VIA 1.518 35.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 35.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.813 1.563 34.847 ;
      VIA 1.518 34.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 34.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 34.273 1.563 34.307 ;
      VIA 1.518 34.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 34.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.733 1.563 33.767 ;
      VIA 1.518 33.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 33.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 33.193 1.563 33.227 ;
      VIA 1.518 33.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 33.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.653 1.563 32.687 ;
      VIA 1.518 32.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 32.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 32.113 1.563 32.147 ;
      VIA 1.518 32.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 32.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.573 1.563 31.607 ;
      VIA 1.518 31.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 31.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 31.033 1.563 31.067 ;
      VIA 1.518 31.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 31.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 30.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 30.493 1.563 30.527 ;
      VIA 1.518 30.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 30.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.953 1.563 29.987 ;
      VIA 1.518 29.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 29.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 29.413 1.563 29.447 ;
      VIA 1.518 29.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 29.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.873 1.563 28.907 ;
      VIA 1.518 28.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 28.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 28.333 1.563 28.367 ;
      VIA 1.518 28.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 28.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.81 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.793 1.563 27.827 ;
      VIA 1.518 27.81 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.81 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 27.27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 27.253 1.563 27.287 ;
      VIA 1.518 27.27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 27.27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.73 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.713 1.563 26.747 ;
      VIA 1.518 26.73 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.73 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 26.19 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 26.173 1.563 26.207 ;
      VIA 1.518 26.19 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 26.19 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.65 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.633 1.563 25.667 ;
      VIA 1.518 25.65 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.65 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 25.11 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 25.093 1.563 25.127 ;
      VIA 1.518 25.11 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 25.11 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.57 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.553 1.563 24.587 ;
      VIA 1.518 24.57 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.57 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 24.03 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 24.013 1.563 24.047 ;
      VIA 1.518 24.03 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 24.03 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 23.49 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 23.473 1.563 23.507 ;
      VIA 1.518 23.49 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 23.49 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.95 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.933 1.563 22.967 ;
      VIA 1.518 22.95 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.95 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 22.41 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 22.393 1.563 22.427 ;
      VIA 1.518 22.41 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 22.41 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.87 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.853 1.563 21.887 ;
      VIA 1.518 21.87 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.87 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 21.33 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 21.313 1.563 21.347 ;
      VIA 1.518 21.33 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 21.33 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.79 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.773 1.563 20.807 ;
      VIA 1.518 20.79 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.79 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 20.25 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 20.233 1.563 20.267 ;
      VIA 1.518 20.25 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 20.25 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.71 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.693 1.563 19.727 ;
      VIA 1.518 19.71 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.71 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 19.17 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 19.153 1.563 19.187 ;
      VIA 1.518 19.17 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 19.17 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.63 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.613 1.563 18.647 ;
      VIA 1.518 18.63 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.63 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 18.09 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 18.073 1.563 18.107 ;
      VIA 1.518 18.09 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 18.09 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.55 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 17.533 1.563 17.567 ;
      VIA 1.518 17.55 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.55 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 17.01 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.993 1.563 17.027 ;
      VIA 1.518 17.01 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 17.01 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 16.47 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 16.453 1.563 16.487 ;
      VIA 1.518 16.47 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 16.47 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.93 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.913 1.563 15.947 ;
      VIA 1.518 15.93 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.93 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 15.39 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 15.373 1.563 15.407 ;
      VIA 1.518 15.39 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 15.39 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.85 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.833 1.563 14.867 ;
      VIA 1.518 14.85 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.85 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 14.31 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 14.293 1.563 14.327 ;
      VIA 1.518 14.31 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 14.31 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.77 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.753 1.563 13.787 ;
      VIA 1.518 13.77 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.77 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 13.23 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 13.213 1.563 13.247 ;
      VIA 1.518 13.23 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 13.23 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.69 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.673 1.563 12.707 ;
      VIA 1.518 12.69 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.69 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 12.15 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 12.133 1.563 12.167 ;
      VIA 1.518 12.15 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 12.15 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.61 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.593 1.563 11.627 ;
      VIA 1.518 11.61 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.61 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 11.07 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.053 1.563 11.087 ;
      VIA 1.518 11.07 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 11.07 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 10.53 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 10.513 1.563 10.547 ;
      VIA 1.518 10.53 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 10.53 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.99 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.973 1.563 10.007 ;
      VIA 1.518 9.99 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.99 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 9.45 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.433 1.563 9.467 ;
      VIA 1.518 9.45 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 9.45 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.91 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.893 1.563 8.927 ;
      VIA 1.518 8.91 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.91 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 8.37 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.353 1.563 8.387 ;
      VIA 1.518 8.37 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 8.37 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.83 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.813 1.563 7.847 ;
      VIA 1.518 7.83 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.83 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 7.29 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.273 1.563 7.307 ;
      VIA 1.518 7.29 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 7.29 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.75 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.733 1.563 6.767 ;
      VIA 1.518 6.75 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.75 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 6.21 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.193 1.563 6.227 ;
      VIA 1.518 6.21 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 6.21 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.67 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.653 1.563 5.687 ;
      VIA 1.518 5.67 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.67 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 5.13 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.113 1.563 5.147 ;
      VIA 1.518 5.13 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 5.13 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.59 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 run_benchmark_VIA23_1_3_36_36 ;
      VIA 20.655 40.23 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 39.69 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 39.15 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 38.61 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 38.07 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 37.53 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 36.99 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 36.45 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 35.91 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 35.37 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 34.83 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 34.29 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 33.75 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 33.21 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 32.67 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 32.13 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 31.59 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 31.05 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 30.51 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 29.97 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 29.43 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 28.89 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 28.35 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 27.81 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 27.27 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 26.73 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 26.19 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 25.65 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 25.11 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 24.57 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 24.03 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 23.49 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 22.95 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 22.41 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 21.87 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 21.33 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 20.79 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 20.25 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 19.71 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 19.17 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 18.63 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 18.09 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 17.55 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 17.01 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 16.47 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 15.93 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 15.39 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 14.85 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 14.31 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 13.77 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 13.23 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 12.69 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 12.15 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 11.61 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 11.07 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 10.53 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 9.99 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 9.45 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 8.91 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 8.37 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 7.83 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 7.29 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 6.75 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 6.21 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 5.67 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 5.13 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 4.59 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 4.05 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 3.51 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 2.97 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 2.43 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 1.89 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 1.35 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.266 37.449 36.81 37.737 ;
        RECT  1.266 31.449 36.81 31.737 ;
        RECT  1.266 25.449 36.81 25.737 ;
        RECT  1.266 19.449 36.81 19.737 ;
        RECT  1.266 13.449 36.81 13.737 ;
        RECT  1.266 7.449 36.81 7.737 ;
        RECT  1.266 1.449 36.81 1.737 ;
      LAYER M5 ;
        RECT  36.69 1.057 36.81 39.983 ;
        RECT  30.786 1.057 30.906 39.983 ;
        RECT  24.882 1.057 25.002 39.983 ;
        RECT  18.978 1.057 19.098 39.983 ;
        RECT  13.074 1.057 13.194 39.983 ;
        RECT  7.17 1.057 7.29 39.983 ;
        RECT  1.266 1.057 1.386 39.983 ;
      LAYER M2 ;
        RECT  1.026 39.951 40.284 39.969 ;
        RECT  1.026 39.411 40.284 39.429 ;
        RECT  1.026 38.871 40.284 38.889 ;
        RECT  1.026 38.331 40.284 38.349 ;
        RECT  1.026 37.791 40.284 37.809 ;
        RECT  1.026 37.251 40.284 37.269 ;
        RECT  1.026 36.711 40.284 36.729 ;
        RECT  1.026 36.171 40.284 36.189 ;
        RECT  1.026 35.631 40.284 35.649 ;
        RECT  1.026 35.091 40.284 35.109 ;
        RECT  1.026 34.551 40.284 34.569 ;
        RECT  1.026 34.011 40.284 34.029 ;
        RECT  1.026 33.471 40.284 33.489 ;
        RECT  1.026 32.931 40.284 32.949 ;
        RECT  1.026 32.391 40.284 32.409 ;
        RECT  1.026 31.851 40.284 31.869 ;
        RECT  1.026 31.311 40.284 31.329 ;
        RECT  1.026 30.771 40.284 30.789 ;
        RECT  1.026 30.231 40.284 30.249 ;
        RECT  1.026 29.691 40.284 29.709 ;
        RECT  1.026 29.151 40.284 29.169 ;
        RECT  1.026 28.611 40.284 28.629 ;
        RECT  1.026 28.071 40.284 28.089 ;
        RECT  1.026 27.531 40.284 27.549 ;
        RECT  1.026 26.991 40.284 27.009 ;
        RECT  1.026 26.451 40.284 26.469 ;
        RECT  1.026 25.911 40.284 25.929 ;
        RECT  1.026 25.371 40.284 25.389 ;
        RECT  1.026 24.831 40.284 24.849 ;
        RECT  1.026 24.291 40.284 24.309 ;
        RECT  1.026 23.751 40.284 23.769 ;
        RECT  1.026 23.211 40.284 23.229 ;
        RECT  1.026 22.671 40.284 22.689 ;
        RECT  1.026 22.131 40.284 22.149 ;
        RECT  1.026 21.591 40.284 21.609 ;
        RECT  1.026 21.051 40.284 21.069 ;
        RECT  1.026 20.511 40.284 20.529 ;
        RECT  1.026 19.971 40.284 19.989 ;
        RECT  1.026 19.431 40.284 19.449 ;
        RECT  1.026 18.891 40.284 18.909 ;
        RECT  1.026 18.351 40.284 18.369 ;
        RECT  1.026 17.811 40.284 17.829 ;
        RECT  1.026 17.271 40.284 17.289 ;
        RECT  1.026 16.731 40.284 16.749 ;
        RECT  1.026 16.191 40.284 16.209 ;
        RECT  1.026 15.651 40.284 15.669 ;
        RECT  1.026 15.111 40.284 15.129 ;
        RECT  1.026 14.571 40.284 14.589 ;
        RECT  1.026 14.031 40.284 14.049 ;
        RECT  1.026 13.491 40.284 13.509 ;
        RECT  1.026 12.951 40.284 12.969 ;
        RECT  1.026 12.411 40.284 12.429 ;
        RECT  1.026 11.871 40.284 11.889 ;
        RECT  1.026 11.331 40.284 11.349 ;
        RECT  1.026 10.791 40.284 10.809 ;
        RECT  1.026 10.251 40.284 10.269 ;
        RECT  1.026 9.711 40.284 9.729 ;
        RECT  1.026 9.171 40.284 9.189 ;
        RECT  1.026 8.631 40.284 8.649 ;
        RECT  1.026 8.091 40.284 8.109 ;
        RECT  1.026 7.551 40.284 7.569 ;
        RECT  1.026 7.011 40.284 7.029 ;
        RECT  1.026 6.471 40.284 6.489 ;
        RECT  1.026 5.931 40.284 5.949 ;
        RECT  1.026 5.391 40.284 5.409 ;
        RECT  1.026 4.851 40.284 4.869 ;
        RECT  1.026 4.311 40.284 4.329 ;
        RECT  1.026 3.771 40.284 3.789 ;
        RECT  1.026 3.231 40.284 3.249 ;
        RECT  1.026 2.691 40.284 2.709 ;
        RECT  1.026 2.151 40.284 2.169 ;
        RECT  1.026 1.611 40.284 1.629 ;
        RECT  1.026 1.071 40.284 1.089 ;
      LAYER M1 ;
        RECT  1.026 39.951 40.284 39.969 ;
        RECT  1.026 39.411 40.284 39.429 ;
        RECT  1.026 38.871 40.284 38.889 ;
        RECT  1.026 38.331 40.284 38.349 ;
        RECT  1.026 37.791 40.284 37.809 ;
        RECT  1.026 37.251 40.284 37.269 ;
        RECT  1.026 36.711 40.284 36.729 ;
        RECT  1.026 36.171 40.284 36.189 ;
        RECT  1.026 35.631 40.284 35.649 ;
        RECT  1.026 35.091 40.284 35.109 ;
        RECT  1.026 34.551 40.284 34.569 ;
        RECT  1.026 34.011 40.284 34.029 ;
        RECT  1.026 33.471 40.284 33.489 ;
        RECT  1.026 32.931 40.284 32.949 ;
        RECT  1.026 32.391 40.284 32.409 ;
        RECT  1.026 31.851 40.284 31.869 ;
        RECT  1.026 31.311 40.284 31.329 ;
        RECT  1.026 30.771 40.284 30.789 ;
        RECT  1.026 30.231 40.284 30.249 ;
        RECT  1.026 29.691 40.284 29.709 ;
        RECT  1.026 29.151 40.284 29.169 ;
        RECT  1.026 28.611 40.284 28.629 ;
        RECT  1.026 28.071 40.284 28.089 ;
        RECT  1.026 27.531 40.284 27.549 ;
        RECT  1.026 26.991 40.284 27.009 ;
        RECT  1.026 26.451 40.284 26.469 ;
        RECT  1.026 25.911 40.284 25.929 ;
        RECT  1.026 25.371 40.284 25.389 ;
        RECT  1.026 24.831 40.284 24.849 ;
        RECT  1.026 24.291 40.284 24.309 ;
        RECT  1.026 23.751 40.284 23.769 ;
        RECT  1.026 23.211 40.284 23.229 ;
        RECT  1.026 22.671 40.284 22.689 ;
        RECT  1.026 22.131 40.284 22.149 ;
        RECT  1.026 21.591 40.284 21.609 ;
        RECT  1.026 21.051 40.284 21.069 ;
        RECT  1.026 20.511 40.284 20.529 ;
        RECT  1.026 19.971 40.284 19.989 ;
        RECT  1.026 19.431 40.284 19.449 ;
        RECT  1.026 18.891 40.284 18.909 ;
        RECT  1.026 18.351 40.284 18.369 ;
        RECT  1.026 17.811 40.284 17.829 ;
        RECT  1.026 17.271 40.284 17.289 ;
        RECT  1.026 16.731 40.284 16.749 ;
        RECT  1.026 16.191 40.284 16.209 ;
        RECT  1.026 15.651 40.284 15.669 ;
        RECT  1.026 15.111 40.284 15.129 ;
        RECT  1.026 14.571 40.284 14.589 ;
        RECT  1.026 14.031 40.284 14.049 ;
        RECT  1.026 13.491 40.284 13.509 ;
        RECT  1.026 12.951 40.284 12.969 ;
        RECT  1.026 12.411 40.284 12.429 ;
        RECT  1.026 11.871 40.284 11.889 ;
        RECT  1.026 11.331 40.284 11.349 ;
        RECT  1.026 10.791 40.284 10.809 ;
        RECT  1.026 10.251 40.284 10.269 ;
        RECT  1.026 9.711 40.284 9.729 ;
        RECT  1.026 9.171 40.284 9.189 ;
        RECT  1.026 8.631 40.284 8.649 ;
        RECT  1.026 8.091 40.284 8.109 ;
        RECT  1.026 7.551 40.284 7.569 ;
        RECT  1.026 7.011 40.284 7.029 ;
        RECT  1.026 6.471 40.284 6.489 ;
        RECT  1.026 5.931 40.284 5.949 ;
        RECT  1.026 5.391 40.284 5.409 ;
        RECT  1.026 4.851 40.284 4.869 ;
        RECT  1.026 4.311 40.284 4.329 ;
        RECT  1.026 3.771 40.284 3.789 ;
        RECT  1.026 3.231 40.284 3.249 ;
        RECT  1.026 2.691 40.284 2.709 ;
        RECT  1.026 2.151 40.284 2.169 ;
        RECT  1.026 1.611 40.284 1.629 ;
        RECT  1.026 1.071 40.284 1.089 ;
      VIA 36.75 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 30.846 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 24.942 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 19.038 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 13.134 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 37.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 31.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 25.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 19.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 13.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 7.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 1.593 run_benchmark_via5_6_120_288_1_2_58_322 ;
      VIA 36.75 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.943 36.795 39.977 ;
      VIA 36.75 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 39.403 36.795 39.437 ;
      VIA 36.75 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.863 36.795 38.897 ;
      VIA 36.75 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 38.323 36.795 38.357 ;
      VIA 36.75 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.783 36.795 37.817 ;
      VIA 36.75 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 37.243 36.795 37.277 ;
      VIA 36.75 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.703 36.795 36.737 ;
      VIA 36.75 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 36.163 36.795 36.197 ;
      VIA 36.75 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.623 36.795 35.657 ;
      VIA 36.75 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 35.083 36.795 35.117 ;
      VIA 36.75 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.543 36.795 34.577 ;
      VIA 36.75 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 34.003 36.795 34.037 ;
      VIA 36.75 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 33.463 36.795 33.497 ;
      VIA 36.75 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.923 36.795 32.957 ;
      VIA 36.75 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 32.383 36.795 32.417 ;
      VIA 36.75 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.843 36.795 31.877 ;
      VIA 36.75 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 31.303 36.795 31.337 ;
      VIA 36.75 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.763 36.795 30.797 ;
      VIA 36.75 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 30.223 36.795 30.257 ;
      VIA 36.75 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.683 36.795 29.717 ;
      VIA 36.75 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 29.143 36.795 29.177 ;
      VIA 36.75 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.603 36.795 28.637 ;
      VIA 36.75 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 28.063 36.795 28.097 ;
      VIA 36.75 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 27.523 36.795 27.557 ;
      VIA 36.75 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.983 36.795 27.017 ;
      VIA 36.75 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 26.443 36.795 26.477 ;
      VIA 36.75 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.903 36.795 25.937 ;
      VIA 36.75 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 25.363 36.795 25.397 ;
      VIA 36.75 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.823 36.795 24.857 ;
      VIA 36.75 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 24.283 36.795 24.317 ;
      VIA 36.75 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.743 36.795 23.777 ;
      VIA 36.75 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 23.203 36.795 23.237 ;
      VIA 36.75 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.663 36.795 22.697 ;
      VIA 36.75 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 22.123 36.795 22.157 ;
      VIA 36.75 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.583 36.795 21.617 ;
      VIA 36.75 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 21.043 36.795 21.077 ;
      VIA 36.75 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 20.503 36.795 20.537 ;
      VIA 36.75 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.963 36.795 19.997 ;
      VIA 36.75 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 19.423 36.795 19.457 ;
      VIA 36.75 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.883 36.795 18.917 ;
      VIA 36.75 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 18.343 36.795 18.377 ;
      VIA 36.75 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.803 36.795 17.837 ;
      VIA 36.75 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 17.263 36.795 17.297 ;
      VIA 36.75 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.723 36.795 16.757 ;
      VIA 36.75 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 16.183 36.795 16.217 ;
      VIA 36.75 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.643 36.795 15.677 ;
      VIA 36.75 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 15.103 36.795 15.137 ;
      VIA 36.75 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.563 36.795 14.597 ;
      VIA 36.75 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 14.023 36.795 14.057 ;
      VIA 36.75 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 13.483 36.795 13.517 ;
      VIA 36.75 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.943 36.795 12.977 ;
      VIA 36.75 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 12.403 36.795 12.437 ;
      VIA 36.75 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.863 36.795 11.897 ;
      VIA 36.75 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 11.323 36.795 11.357 ;
      VIA 36.75 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.783 36.795 10.817 ;
      VIA 36.75 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 10.243 36.795 10.277 ;
      VIA 36.75 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.703 36.795 9.737 ;
      VIA 36.75 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 9.163 36.795 9.197 ;
      VIA 36.75 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.623 36.795 8.657 ;
      VIA 36.75 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 8.083 36.795 8.117 ;
      VIA 36.75 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.543 36.795 7.577 ;
      VIA 36.75 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 7.003 36.795 7.037 ;
      VIA 36.75 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 6.463 36.795 6.497 ;
      VIA 36.75 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.923 36.795 5.957 ;
      VIA 36.75 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 5.383 36.795 5.417 ;
      VIA 36.75 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.843 36.795 4.877 ;
      VIA 36.75 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 4.303 36.795 4.337 ;
      VIA 36.75 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.763 36.795 3.797 ;
      VIA 36.75 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 3.223 36.795 3.257 ;
      VIA 36.75 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.683 36.795 2.717 ;
      VIA 36.75 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 2.143 36.795 2.177 ;
      VIA 36.75 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.603 36.795 1.637 ;
      VIA 36.75 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 36.75 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  36.705 1.063 36.795 1.097 ;
      VIA 36.75 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 36.75 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.943 30.891 39.977 ;
      VIA 30.846 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 39.403 30.891 39.437 ;
      VIA 30.846 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.863 30.891 38.897 ;
      VIA 30.846 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 38.323 30.891 38.357 ;
      VIA 30.846 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.783 30.891 37.817 ;
      VIA 30.846 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 37.243 30.891 37.277 ;
      VIA 30.846 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.703 30.891 36.737 ;
      VIA 30.846 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 36.163 30.891 36.197 ;
      VIA 30.846 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.623 30.891 35.657 ;
      VIA 30.846 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 35.083 30.891 35.117 ;
      VIA 30.846 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.543 30.891 34.577 ;
      VIA 30.846 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 34.003 30.891 34.037 ;
      VIA 30.846 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 33.463 30.891 33.497 ;
      VIA 30.846 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.923 30.891 32.957 ;
      VIA 30.846 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 32.383 30.891 32.417 ;
      VIA 30.846 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.843 30.891 31.877 ;
      VIA 30.846 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 31.303 30.891 31.337 ;
      VIA 30.846 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.763 30.891 30.797 ;
      VIA 30.846 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 30.223 30.891 30.257 ;
      VIA 30.846 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.683 30.891 29.717 ;
      VIA 30.846 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 29.143 30.891 29.177 ;
      VIA 30.846 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.603 30.891 28.637 ;
      VIA 30.846 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 28.063 30.891 28.097 ;
      VIA 30.846 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 27.523 30.891 27.557 ;
      VIA 30.846 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.983 30.891 27.017 ;
      VIA 30.846 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 26.443 30.891 26.477 ;
      VIA 30.846 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.903 30.891 25.937 ;
      VIA 30.846 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 25.363 30.891 25.397 ;
      VIA 30.846 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.823 30.891 24.857 ;
      VIA 30.846 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 24.283 30.891 24.317 ;
      VIA 30.846 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.743 30.891 23.777 ;
      VIA 30.846 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 23.203 30.891 23.237 ;
      VIA 30.846 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.663 30.891 22.697 ;
      VIA 30.846 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 22.123 30.891 22.157 ;
      VIA 30.846 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.583 30.891 21.617 ;
      VIA 30.846 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 21.043 30.891 21.077 ;
      VIA 30.846 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 20.503 30.891 20.537 ;
      VIA 30.846 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.963 30.891 19.997 ;
      VIA 30.846 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 19.423 30.891 19.457 ;
      VIA 30.846 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.883 30.891 18.917 ;
      VIA 30.846 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 18.343 30.891 18.377 ;
      VIA 30.846 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.803 30.891 17.837 ;
      VIA 30.846 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 17.263 30.891 17.297 ;
      VIA 30.846 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.723 30.891 16.757 ;
      VIA 30.846 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 16.183 30.891 16.217 ;
      VIA 30.846 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.643 30.891 15.677 ;
      VIA 30.846 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 15.103 30.891 15.137 ;
      VIA 30.846 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.563 30.891 14.597 ;
      VIA 30.846 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 14.023 30.891 14.057 ;
      VIA 30.846 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 13.483 30.891 13.517 ;
      VIA 30.846 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.943 30.891 12.977 ;
      VIA 30.846 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 12.403 30.891 12.437 ;
      VIA 30.846 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.863 30.891 11.897 ;
      VIA 30.846 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 11.323 30.891 11.357 ;
      VIA 30.846 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.783 30.891 10.817 ;
      VIA 30.846 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 10.243 30.891 10.277 ;
      VIA 30.846 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.703 30.891 9.737 ;
      VIA 30.846 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 9.163 30.891 9.197 ;
      VIA 30.846 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.623 30.891 8.657 ;
      VIA 30.846 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 8.083 30.891 8.117 ;
      VIA 30.846 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.543 30.891 7.577 ;
      VIA 30.846 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 7.003 30.891 7.037 ;
      VIA 30.846 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 6.463 30.891 6.497 ;
      VIA 30.846 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.923 30.891 5.957 ;
      VIA 30.846 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 5.383 30.891 5.417 ;
      VIA 30.846 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.843 30.891 4.877 ;
      VIA 30.846 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 4.303 30.891 4.337 ;
      VIA 30.846 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.763 30.891 3.797 ;
      VIA 30.846 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 3.223 30.891 3.257 ;
      VIA 30.846 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.683 30.891 2.717 ;
      VIA 30.846 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 2.143 30.891 2.177 ;
      VIA 30.846 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.603 30.891 1.637 ;
      VIA 30.846 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 30.846 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  30.801 1.063 30.891 1.097 ;
      VIA 30.846 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 30.846 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.943 24.987 39.977 ;
      VIA 24.942 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 39.403 24.987 39.437 ;
      VIA 24.942 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.863 24.987 38.897 ;
      VIA 24.942 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 38.323 24.987 38.357 ;
      VIA 24.942 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.783 24.987 37.817 ;
      VIA 24.942 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 37.243 24.987 37.277 ;
      VIA 24.942 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.703 24.987 36.737 ;
      VIA 24.942 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 36.163 24.987 36.197 ;
      VIA 24.942 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.623 24.987 35.657 ;
      VIA 24.942 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 35.083 24.987 35.117 ;
      VIA 24.942 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.543 24.987 34.577 ;
      VIA 24.942 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 34.003 24.987 34.037 ;
      VIA 24.942 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 33.463 24.987 33.497 ;
      VIA 24.942 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.923 24.987 32.957 ;
      VIA 24.942 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 32.383 24.987 32.417 ;
      VIA 24.942 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.843 24.987 31.877 ;
      VIA 24.942 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 31.303 24.987 31.337 ;
      VIA 24.942 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.763 24.987 30.797 ;
      VIA 24.942 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 30.223 24.987 30.257 ;
      VIA 24.942 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.683 24.987 29.717 ;
      VIA 24.942 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 29.143 24.987 29.177 ;
      VIA 24.942 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.603 24.987 28.637 ;
      VIA 24.942 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 28.063 24.987 28.097 ;
      VIA 24.942 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 27.523 24.987 27.557 ;
      VIA 24.942 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.983 24.987 27.017 ;
      VIA 24.942 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 26.443 24.987 26.477 ;
      VIA 24.942 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.903 24.987 25.937 ;
      VIA 24.942 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 25.363 24.987 25.397 ;
      VIA 24.942 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.823 24.987 24.857 ;
      VIA 24.942 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 24.283 24.987 24.317 ;
      VIA 24.942 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.743 24.987 23.777 ;
      VIA 24.942 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 23.203 24.987 23.237 ;
      VIA 24.942 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.663 24.987 22.697 ;
      VIA 24.942 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 22.123 24.987 22.157 ;
      VIA 24.942 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.583 24.987 21.617 ;
      VIA 24.942 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 21.043 24.987 21.077 ;
      VIA 24.942 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 20.503 24.987 20.537 ;
      VIA 24.942 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.963 24.987 19.997 ;
      VIA 24.942 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 19.423 24.987 19.457 ;
      VIA 24.942 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.883 24.987 18.917 ;
      VIA 24.942 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 18.343 24.987 18.377 ;
      VIA 24.942 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.803 24.987 17.837 ;
      VIA 24.942 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 17.263 24.987 17.297 ;
      VIA 24.942 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.723 24.987 16.757 ;
      VIA 24.942 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 16.183 24.987 16.217 ;
      VIA 24.942 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.643 24.987 15.677 ;
      VIA 24.942 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 15.103 24.987 15.137 ;
      VIA 24.942 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.563 24.987 14.597 ;
      VIA 24.942 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 14.023 24.987 14.057 ;
      VIA 24.942 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 13.483 24.987 13.517 ;
      VIA 24.942 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.943 24.987 12.977 ;
      VIA 24.942 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 12.403 24.987 12.437 ;
      VIA 24.942 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.863 24.987 11.897 ;
      VIA 24.942 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 11.323 24.987 11.357 ;
      VIA 24.942 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.783 24.987 10.817 ;
      VIA 24.942 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 10.243 24.987 10.277 ;
      VIA 24.942 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.703 24.987 9.737 ;
      VIA 24.942 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 9.163 24.987 9.197 ;
      VIA 24.942 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.623 24.987 8.657 ;
      VIA 24.942 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 8.083 24.987 8.117 ;
      VIA 24.942 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.543 24.987 7.577 ;
      VIA 24.942 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 7.003 24.987 7.037 ;
      VIA 24.942 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 6.463 24.987 6.497 ;
      VIA 24.942 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.923 24.987 5.957 ;
      VIA 24.942 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 5.383 24.987 5.417 ;
      VIA 24.942 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.843 24.987 4.877 ;
      VIA 24.942 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 4.303 24.987 4.337 ;
      VIA 24.942 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.763 24.987 3.797 ;
      VIA 24.942 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 3.223 24.987 3.257 ;
      VIA 24.942 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.683 24.987 2.717 ;
      VIA 24.942 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 2.143 24.987 2.177 ;
      VIA 24.942 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.603 24.987 1.637 ;
      VIA 24.942 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 24.942 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  24.897 1.063 24.987 1.097 ;
      VIA 24.942 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 24.942 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.943 19.083 39.977 ;
      VIA 19.038 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 39.403 19.083 39.437 ;
      VIA 19.038 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.863 19.083 38.897 ;
      VIA 19.038 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 38.323 19.083 38.357 ;
      VIA 19.038 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.783 19.083 37.817 ;
      VIA 19.038 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 37.243 19.083 37.277 ;
      VIA 19.038 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.703 19.083 36.737 ;
      VIA 19.038 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 36.163 19.083 36.197 ;
      VIA 19.038 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.623 19.083 35.657 ;
      VIA 19.038 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 35.083 19.083 35.117 ;
      VIA 19.038 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.543 19.083 34.577 ;
      VIA 19.038 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 34.003 19.083 34.037 ;
      VIA 19.038 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 33.463 19.083 33.497 ;
      VIA 19.038 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.923 19.083 32.957 ;
      VIA 19.038 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 32.383 19.083 32.417 ;
      VIA 19.038 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.843 19.083 31.877 ;
      VIA 19.038 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 31.303 19.083 31.337 ;
      VIA 19.038 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.763 19.083 30.797 ;
      VIA 19.038 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 30.223 19.083 30.257 ;
      VIA 19.038 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.683 19.083 29.717 ;
      VIA 19.038 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 29.143 19.083 29.177 ;
      VIA 19.038 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.603 19.083 28.637 ;
      VIA 19.038 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 28.063 19.083 28.097 ;
      VIA 19.038 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 27.523 19.083 27.557 ;
      VIA 19.038 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.983 19.083 27.017 ;
      VIA 19.038 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 26.443 19.083 26.477 ;
      VIA 19.038 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.903 19.083 25.937 ;
      VIA 19.038 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 25.363 19.083 25.397 ;
      VIA 19.038 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.823 19.083 24.857 ;
      VIA 19.038 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 24.283 19.083 24.317 ;
      VIA 19.038 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.743 19.083 23.777 ;
      VIA 19.038 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 23.203 19.083 23.237 ;
      VIA 19.038 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.663 19.083 22.697 ;
      VIA 19.038 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 22.123 19.083 22.157 ;
      VIA 19.038 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.583 19.083 21.617 ;
      VIA 19.038 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 21.043 19.083 21.077 ;
      VIA 19.038 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 20.503 19.083 20.537 ;
      VIA 19.038 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.963 19.083 19.997 ;
      VIA 19.038 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 19.423 19.083 19.457 ;
      VIA 19.038 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.883 19.083 18.917 ;
      VIA 19.038 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 18.343 19.083 18.377 ;
      VIA 19.038 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.803 19.083 17.837 ;
      VIA 19.038 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 17.263 19.083 17.297 ;
      VIA 19.038 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.723 19.083 16.757 ;
      VIA 19.038 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 16.183 19.083 16.217 ;
      VIA 19.038 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.643 19.083 15.677 ;
      VIA 19.038 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 15.103 19.083 15.137 ;
      VIA 19.038 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.563 19.083 14.597 ;
      VIA 19.038 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 14.023 19.083 14.057 ;
      VIA 19.038 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 13.483 19.083 13.517 ;
      VIA 19.038 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.943 19.083 12.977 ;
      VIA 19.038 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 12.403 19.083 12.437 ;
      VIA 19.038 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.863 19.083 11.897 ;
      VIA 19.038 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 11.323 19.083 11.357 ;
      VIA 19.038 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.783 19.083 10.817 ;
      VIA 19.038 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 10.243 19.083 10.277 ;
      VIA 19.038 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.703 19.083 9.737 ;
      VIA 19.038 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 9.163 19.083 9.197 ;
      VIA 19.038 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.623 19.083 8.657 ;
      VIA 19.038 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 8.083 19.083 8.117 ;
      VIA 19.038 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.543 19.083 7.577 ;
      VIA 19.038 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 7.003 19.083 7.037 ;
      VIA 19.038 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 6.463 19.083 6.497 ;
      VIA 19.038 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.923 19.083 5.957 ;
      VIA 19.038 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 5.383 19.083 5.417 ;
      VIA 19.038 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.843 19.083 4.877 ;
      VIA 19.038 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 4.303 19.083 4.337 ;
      VIA 19.038 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.763 19.083 3.797 ;
      VIA 19.038 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 3.223 19.083 3.257 ;
      VIA 19.038 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.683 19.083 2.717 ;
      VIA 19.038 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 2.143 19.083 2.177 ;
      VIA 19.038 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.603 19.083 1.637 ;
      VIA 19.038 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 19.038 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  18.993 1.063 19.083 1.097 ;
      VIA 19.038 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 19.038 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.943 13.179 39.977 ;
      VIA 13.134 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 39.403 13.179 39.437 ;
      VIA 13.134 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.863 13.179 38.897 ;
      VIA 13.134 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 38.323 13.179 38.357 ;
      VIA 13.134 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.783 13.179 37.817 ;
      VIA 13.134 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 37.243 13.179 37.277 ;
      VIA 13.134 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.703 13.179 36.737 ;
      VIA 13.134 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 36.163 13.179 36.197 ;
      VIA 13.134 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.623 13.179 35.657 ;
      VIA 13.134 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 35.083 13.179 35.117 ;
      VIA 13.134 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.543 13.179 34.577 ;
      VIA 13.134 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 34.003 13.179 34.037 ;
      VIA 13.134 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 33.463 13.179 33.497 ;
      VIA 13.134 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.923 13.179 32.957 ;
      VIA 13.134 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 32.383 13.179 32.417 ;
      VIA 13.134 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.843 13.179 31.877 ;
      VIA 13.134 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 31.303 13.179 31.337 ;
      VIA 13.134 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.763 13.179 30.797 ;
      VIA 13.134 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 30.223 13.179 30.257 ;
      VIA 13.134 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.683 13.179 29.717 ;
      VIA 13.134 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 29.143 13.179 29.177 ;
      VIA 13.134 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.603 13.179 28.637 ;
      VIA 13.134 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 28.063 13.179 28.097 ;
      VIA 13.134 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 27.523 13.179 27.557 ;
      VIA 13.134 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.983 13.179 27.017 ;
      VIA 13.134 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 26.443 13.179 26.477 ;
      VIA 13.134 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.903 13.179 25.937 ;
      VIA 13.134 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 25.363 13.179 25.397 ;
      VIA 13.134 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.823 13.179 24.857 ;
      VIA 13.134 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 24.283 13.179 24.317 ;
      VIA 13.134 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.743 13.179 23.777 ;
      VIA 13.134 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 23.203 13.179 23.237 ;
      VIA 13.134 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.663 13.179 22.697 ;
      VIA 13.134 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 22.123 13.179 22.157 ;
      VIA 13.134 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.583 13.179 21.617 ;
      VIA 13.134 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 21.043 13.179 21.077 ;
      VIA 13.134 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 20.503 13.179 20.537 ;
      VIA 13.134 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.963 13.179 19.997 ;
      VIA 13.134 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 19.423 13.179 19.457 ;
      VIA 13.134 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.883 13.179 18.917 ;
      VIA 13.134 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 18.343 13.179 18.377 ;
      VIA 13.134 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.803 13.179 17.837 ;
      VIA 13.134 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 17.263 13.179 17.297 ;
      VIA 13.134 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.723 13.179 16.757 ;
      VIA 13.134 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 16.183 13.179 16.217 ;
      VIA 13.134 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.643 13.179 15.677 ;
      VIA 13.134 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 15.103 13.179 15.137 ;
      VIA 13.134 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.563 13.179 14.597 ;
      VIA 13.134 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 14.023 13.179 14.057 ;
      VIA 13.134 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 13.483 13.179 13.517 ;
      VIA 13.134 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.943 13.179 12.977 ;
      VIA 13.134 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 12.403 13.179 12.437 ;
      VIA 13.134 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.863 13.179 11.897 ;
      VIA 13.134 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 11.323 13.179 11.357 ;
      VIA 13.134 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.783 13.179 10.817 ;
      VIA 13.134 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 10.243 13.179 10.277 ;
      VIA 13.134 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.703 13.179 9.737 ;
      VIA 13.134 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 9.163 13.179 9.197 ;
      VIA 13.134 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.623 13.179 8.657 ;
      VIA 13.134 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 8.083 13.179 8.117 ;
      VIA 13.134 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.543 13.179 7.577 ;
      VIA 13.134 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 7.003 13.179 7.037 ;
      VIA 13.134 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 6.463 13.179 6.497 ;
      VIA 13.134 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.923 13.179 5.957 ;
      VIA 13.134 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 5.383 13.179 5.417 ;
      VIA 13.134 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.843 13.179 4.877 ;
      VIA 13.134 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 4.303 13.179 4.337 ;
      VIA 13.134 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.763 13.179 3.797 ;
      VIA 13.134 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 3.223 13.179 3.257 ;
      VIA 13.134 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.683 13.179 2.717 ;
      VIA 13.134 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 2.143 13.179 2.177 ;
      VIA 13.134 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.603 13.179 1.637 ;
      VIA 13.134 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 13.134 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  13.089 1.063 13.179 1.097 ;
      VIA 13.134 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 13.134 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.943 7.275 39.977 ;
      VIA 7.23 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 39.403 7.275 39.437 ;
      VIA 7.23 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.863 7.275 38.897 ;
      VIA 7.23 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 38.323 7.275 38.357 ;
      VIA 7.23 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.783 7.275 37.817 ;
      VIA 7.23 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 37.243 7.275 37.277 ;
      VIA 7.23 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.703 7.275 36.737 ;
      VIA 7.23 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 36.163 7.275 36.197 ;
      VIA 7.23 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.623 7.275 35.657 ;
      VIA 7.23 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 35.083 7.275 35.117 ;
      VIA 7.23 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.543 7.275 34.577 ;
      VIA 7.23 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 34.003 7.275 34.037 ;
      VIA 7.23 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 33.463 7.275 33.497 ;
      VIA 7.23 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.923 7.275 32.957 ;
      VIA 7.23 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 32.383 7.275 32.417 ;
      VIA 7.23 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.843 7.275 31.877 ;
      VIA 7.23 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 31.303 7.275 31.337 ;
      VIA 7.23 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.763 7.275 30.797 ;
      VIA 7.23 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 30.223 7.275 30.257 ;
      VIA 7.23 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.683 7.275 29.717 ;
      VIA 7.23 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 29.143 7.275 29.177 ;
      VIA 7.23 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.603 7.275 28.637 ;
      VIA 7.23 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 28.063 7.275 28.097 ;
      VIA 7.23 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 27.523 7.275 27.557 ;
      VIA 7.23 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.983 7.275 27.017 ;
      VIA 7.23 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 26.443 7.275 26.477 ;
      VIA 7.23 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.903 7.275 25.937 ;
      VIA 7.23 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 25.363 7.275 25.397 ;
      VIA 7.23 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.823 7.275 24.857 ;
      VIA 7.23 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 24.283 7.275 24.317 ;
      VIA 7.23 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.743 7.275 23.777 ;
      VIA 7.23 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 23.203 7.275 23.237 ;
      VIA 7.23 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.663 7.275 22.697 ;
      VIA 7.23 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 22.123 7.275 22.157 ;
      VIA 7.23 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.583 7.275 21.617 ;
      VIA 7.23 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 21.043 7.275 21.077 ;
      VIA 7.23 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 20.503 7.275 20.537 ;
      VIA 7.23 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.963 7.275 19.997 ;
      VIA 7.23 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 19.423 7.275 19.457 ;
      VIA 7.23 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.883 7.275 18.917 ;
      VIA 7.23 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 18.343 7.275 18.377 ;
      VIA 7.23 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.803 7.275 17.837 ;
      VIA 7.23 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 17.263 7.275 17.297 ;
      VIA 7.23 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.723 7.275 16.757 ;
      VIA 7.23 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 16.183 7.275 16.217 ;
      VIA 7.23 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.643 7.275 15.677 ;
      VIA 7.23 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 15.103 7.275 15.137 ;
      VIA 7.23 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.563 7.275 14.597 ;
      VIA 7.23 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 14.023 7.275 14.057 ;
      VIA 7.23 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 13.483 7.275 13.517 ;
      VIA 7.23 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.943 7.275 12.977 ;
      VIA 7.23 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 12.403 7.275 12.437 ;
      VIA 7.23 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.863 7.275 11.897 ;
      VIA 7.23 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.323 7.275 11.357 ;
      VIA 7.23 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.783 7.275 10.817 ;
      VIA 7.23 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.243 7.275 10.277 ;
      VIA 7.23 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.703 7.275 9.737 ;
      VIA 7.23 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.163 7.275 9.197 ;
      VIA 7.23 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.623 7.275 8.657 ;
      VIA 7.23 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.083 7.275 8.117 ;
      VIA 7.23 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.543 7.275 7.577 ;
      VIA 7.23 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.003 7.275 7.037 ;
      VIA 7.23 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 6.463 7.275 6.497 ;
      VIA 7.23 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.923 7.275 5.957 ;
      VIA 7.23 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.383 7.275 5.417 ;
      VIA 7.23 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.843 7.275 4.877 ;
      VIA 7.23 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.303 7.275 4.337 ;
      VIA 7.23 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.763 7.275 3.797 ;
      VIA 7.23 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.223 7.275 3.257 ;
      VIA 7.23 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.683 7.275 2.717 ;
      VIA 7.23 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.143 7.275 2.177 ;
      VIA 7.23 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.603 7.275 1.637 ;
      VIA 7.23 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 7.23 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.063 7.275 1.097 ;
      VIA 7.23 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 7.23 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.943 1.371 39.977 ;
      VIA 1.326 39.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 39.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 39.403 1.371 39.437 ;
      VIA 1.326 39.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 39.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.863 1.371 38.897 ;
      VIA 1.326 38.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 38.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 38.323 1.371 38.357 ;
      VIA 1.326 38.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 38.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.783 1.371 37.817 ;
      VIA 1.326 37.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 37.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 37.243 1.371 37.277 ;
      VIA 1.326 37.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 37.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.703 1.371 36.737 ;
      VIA 1.326 36.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 36.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 36.163 1.371 36.197 ;
      VIA 1.326 36.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 36.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.623 1.371 35.657 ;
      VIA 1.326 35.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 35.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 35.083 1.371 35.117 ;
      VIA 1.326 35.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 35.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.543 1.371 34.577 ;
      VIA 1.326 34.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 34.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 34.003 1.371 34.037 ;
      VIA 1.326 34.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 34.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 33.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 33.463 1.371 33.497 ;
      VIA 1.326 33.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 33.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.923 1.371 32.957 ;
      VIA 1.326 32.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 32.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 32.383 1.371 32.417 ;
      VIA 1.326 32.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 32.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.843 1.371 31.877 ;
      VIA 1.326 31.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 31.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 31.303 1.371 31.337 ;
      VIA 1.326 31.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 31.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.763 1.371 30.797 ;
      VIA 1.326 30.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 30.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 30.223 1.371 30.257 ;
      VIA 1.326 30.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 30.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.683 1.371 29.717 ;
      VIA 1.326 29.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 29.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 29.143 1.371 29.177 ;
      VIA 1.326 29.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 29.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.603 1.371 28.637 ;
      VIA 1.326 28.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 28.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 28.063 1.371 28.097 ;
      VIA 1.326 28.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 28.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27.54 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 27.523 1.371 27.557 ;
      VIA 1.326 27.54 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27.54 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 27 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.983 1.371 27.017 ;
      VIA 1.326 27 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 27 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 26.46 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 26.443 1.371 26.477 ;
      VIA 1.326 26.46 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 26.46 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.92 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.903 1.371 25.937 ;
      VIA 1.326 25.92 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.92 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 25.38 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 25.363 1.371 25.397 ;
      VIA 1.326 25.38 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 25.38 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.84 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.823 1.371 24.857 ;
      VIA 1.326 24.84 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.84 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 24.3 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 24.283 1.371 24.317 ;
      VIA 1.326 24.3 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 24.3 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.76 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.743 1.371 23.777 ;
      VIA 1.326 23.76 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.76 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 23.22 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 23.203 1.371 23.237 ;
      VIA 1.326 23.22 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 23.22 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.68 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.663 1.371 22.697 ;
      VIA 1.326 22.68 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.68 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 22.14 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 22.123 1.371 22.157 ;
      VIA 1.326 22.14 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 22.14 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.6 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.583 1.371 21.617 ;
      VIA 1.326 21.6 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.6 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 21.06 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 21.043 1.371 21.077 ;
      VIA 1.326 21.06 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 21.06 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 20.52 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 20.503 1.371 20.537 ;
      VIA 1.326 20.52 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 20.52 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.98 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.963 1.371 19.997 ;
      VIA 1.326 19.98 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.98 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 19.44 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 19.423 1.371 19.457 ;
      VIA 1.326 19.44 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 19.44 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.9 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.883 1.371 18.917 ;
      VIA 1.326 18.9 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.9 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 18.36 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 18.343 1.371 18.377 ;
      VIA 1.326 18.36 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 18.36 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.82 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.803 1.371 17.837 ;
      VIA 1.326 17.82 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.82 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 17.28 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 17.263 1.371 17.297 ;
      VIA 1.326 17.28 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 17.28 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.74 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.723 1.371 16.757 ;
      VIA 1.326 16.74 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.74 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 16.2 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 16.183 1.371 16.217 ;
      VIA 1.326 16.2 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 16.2 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.66 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.643 1.371 15.677 ;
      VIA 1.326 15.66 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.66 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 15.12 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 15.103 1.371 15.137 ;
      VIA 1.326 15.12 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 15.12 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.58 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.563 1.371 14.597 ;
      VIA 1.326 14.58 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.58 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 14.04 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 14.023 1.371 14.057 ;
      VIA 1.326 14.04 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 14.04 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 13.5 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 13.483 1.371 13.517 ;
      VIA 1.326 13.5 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 13.5 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.96 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.943 1.371 12.977 ;
      VIA 1.326 12.96 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.96 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 12.42 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 12.403 1.371 12.437 ;
      VIA 1.326 12.42 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 12.42 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.88 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.863 1.371 11.897 ;
      VIA 1.326 11.88 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.88 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 11.34 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.323 1.371 11.357 ;
      VIA 1.326 11.34 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 11.34 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.8 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.783 1.371 10.817 ;
      VIA 1.326 10.8 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.8 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 10.26 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.243 1.371 10.277 ;
      VIA 1.326 10.26 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 10.26 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.72 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.703 1.371 9.737 ;
      VIA 1.326 9.72 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.72 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 9.18 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.163 1.371 9.197 ;
      VIA 1.326 9.18 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 9.18 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.64 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.623 1.371 8.657 ;
      VIA 1.326 8.64 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.64 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 8.1 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.083 1.371 8.117 ;
      VIA 1.326 8.1 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 8.1 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.56 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.543 1.371 7.577 ;
      VIA 1.326 7.56 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.56 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 7.02 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.003 1.371 7.037 ;
      VIA 1.326 7.02 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 7.02 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 6.48 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 6.463 1.371 6.497 ;
      VIA 1.326 6.48 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 6.48 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.94 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.923 1.371 5.957 ;
      VIA 1.326 5.94 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.94 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 5.4 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.383 1.371 5.417 ;
      VIA 1.326 5.4 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 5.4 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.86 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 run_benchmark_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 run_benchmark_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 run_benchmark_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 run_benchmark_VIA23_1_3_36_36 ;
      VIA 20.655 39.96 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 39.42 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 38.88 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 38.34 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 37.8 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 37.26 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 36.72 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 36.18 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 35.64 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 35.1 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 34.56 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 34.02 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 33.48 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 32.94 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 32.4 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 31.86 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 31.32 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 30.78 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 30.24 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 29.7 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 29.16 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 28.62 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 28.08 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 27.54 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 27 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 26.46 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 25.92 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 25.38 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 24.84 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 24.3 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 23.76 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 23.22 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 22.68 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 22.14 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 21.6 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 21.06 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 20.52 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 19.98 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 19.44 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 18.9 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 18.36 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 17.82 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 17.28 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 16.74 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 16.2 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 15.66 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 15.12 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 14.58 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 14.04 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 13.5 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 12.96 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 12.42 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 11.88 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 11.34 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 10.8 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 10.26 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 9.72 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 9.18 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 8.64 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 8.1 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 7.56 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 7.02 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 6.48 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 5.94 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 5.4 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 4.86 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 4.32 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 3.78 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 3.24 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 2.7 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 2.16 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 1.62 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
      VIA 20.655 1.08 run_benchmark_via1_2_39258_18_1_1090_36_36 ;
    END
  END VSS
  PIN M_DataRdy[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.672 0 0.696 0.084 ;
    END
  END M_DataRdy[0]
  PIN M_DataRdy[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.768 0 0.792 0.084 ;
    END
  END M_DataRdy[1]
  PIN M_Rdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.984 41.235 10.008 41.319 ;
    END
  END M_Rdata_ram[0]
  PIN M_Rdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.696 0.084 21.72 ;
    END
  END M_Rdata_ram[10]
  PIN M_Rdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.064 0.084 20.088 ;
    END
  END M_Rdata_ram[11]
  PIN M_Rdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.624 0.084 18.648 ;
    END
  END M_Rdata_ram[12]
  PIN M_Rdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.28 0.084 17.304 ;
    END
  END M_Rdata_ram[13]
  PIN M_Rdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.088 0.084 17.112 ;
    END
  END M_Rdata_ram[14]
  PIN M_Rdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.896 0.084 16.92 ;
    END
  END M_Rdata_ram[15]
  PIN M_Rdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.096 0.084 12.12 ;
    END
  END M_Rdata_ram[16]
  PIN M_Rdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.752 0.084 10.776 ;
    END
  END M_Rdata_ram[17]
  PIN M_Rdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.352 0 8.376 0.084 ;
    END
  END M_Rdata_ram[18]
  PIN M_Rdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.448 0 8.472 0.084 ;
    END
  END M_Rdata_ram[19]
  PIN M_Rdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.464 41.235 10.488 41.319 ;
    END
  END M_Rdata_ram[1]
  PIN M_Rdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.544 0 8.568 0.084 ;
    END
  END M_Rdata_ram[20]
  PIN M_Rdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.248 0.084 13.272 ;
    END
  END M_Rdata_ram[21]
  PIN M_Rdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.712 0.084 11.736 ;
    END
  END M_Rdata_ram[22]
  PIN M_Rdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.576 0.084 12.6 ;
    END
  END M_Rdata_ram[23]
  PIN M_Rdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.56 0.084 10.584 ;
    END
  END M_Rdata_ram[24]
  PIN M_Rdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.656 0.084 10.68 ;
    END
  END M_Rdata_ram[25]
  PIN M_Rdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.808 0.084 11.832 ;
    END
  END M_Rdata_ram[26]
  PIN M_Rdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.904 0.084 11.928 ;
    END
  END M_Rdata_ram[27]
  PIN M_Rdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.48 0.084 12.504 ;
    END
  END M_Rdata_ram[28]
  PIN M_Rdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.536 0.084 13.56 ;
    END
  END M_Rdata_ram[29]
  PIN M_Rdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.08 41.235 10.104 41.319 ;
    END
  END M_Rdata_ram[2]
  PIN M_Rdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.496 0.084 14.52 ;
    END
  END M_Rdata_ram[30]
  PIN M_Rdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 32.64 0.084 32.664 ;
    END
  END M_Rdata_ram[31]
  PIN M_Rdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.4 41.235 14.424 41.319 ;
    END
  END M_Rdata_ram[32]
  PIN M_Rdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.304 41.235 14.328 41.319 ;
    END
  END M_Rdata_ram[33]
  PIN M_Rdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.728 41.235 13.752 41.319 ;
    END
  END M_Rdata_ram[34]
  PIN M_Rdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.92 41.235 13.944 41.319 ;
    END
  END M_Rdata_ram[35]
  PIN M_Rdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.208 41.235 14.232 41.319 ;
    END
  END M_Rdata_ram[36]
  PIN M_Rdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.496 41.235 14.52 41.319 ;
    END
  END M_Rdata_ram[37]
  PIN M_Rdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.824 41.235 13.848 41.319 ;
    END
  END M_Rdata_ram[38]
  PIN M_Rdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.016 41.235 14.04 41.319 ;
    END
  END M_Rdata_ram[39]
  PIN M_Rdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 36.192 0.084 36.216 ;
    END
  END M_Rdata_ram[3]
  PIN M_Rdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.112 41.235 14.136 41.319 ;
    END
  END M_Rdata_ram[40]
  PIN M_Rdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.408 0.084 21.432 ;
    END
  END M_Rdata_ram[41]
  PIN M_Rdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.024 0.084 21.048 ;
    END
  END M_Rdata_ram[42]
  PIN M_Rdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.488 0.084 19.512 ;
    END
  END M_Rdata_ram[43]
  PIN M_Rdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.336 0.084 18.36 ;
    END
  END M_Rdata_ram[44]
  PIN M_Rdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.184 0.084 17.208 ;
    END
  END M_Rdata_ram[45]
  PIN M_Rdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.8 0.084 16.824 ;
    END
  END M_Rdata_ram[46]
  PIN M_Rdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.72 0.084 18.744 ;
    END
  END M_Rdata_ram[47]
  PIN M_Rdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.152 0.084 13.176 ;
    END
  END M_Rdata_ram[48]
  PIN M_Rdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.416 0 16.44 0.084 ;
    END
  END M_Rdata_ram[49]
  PIN M_Rdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.272 41.235 10.296 41.319 ;
    END
  END M_Rdata_ram[4]
  PIN M_Rdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.128 0 16.152 0.084 ;
    END
  END M_Rdata_ram[50]
  PIN M_Rdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.208 0 14.232 0.084 ;
    END
  END M_Rdata_ram[51]
  PIN M_Rdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.96 0 12.984 0.084 ;
    END
  END M_Rdata_ram[52]
  PIN M_Rdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.616 0 11.64 0.084 ;
    END
  END M_Rdata_ram[53]
  PIN M_Rdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.096 0 12.12 0.084 ;
    END
  END M_Rdata_ram[54]
  PIN M_Rdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.688 0.084 14.712 ;
    END
  END M_Rdata_ram[55]
  PIN M_Rdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.056 0.084 13.08 ;
    END
  END M_Rdata_ram[56]
  PIN M_Rdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.632 0.084 13.656 ;
    END
  END M_Rdata_ram[57]
  PIN M_Rdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.512 0.084 16.536 ;
    END
  END M_Rdata_ram[58]
  PIN M_Rdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.992 0.084 17.016 ;
    END
  END M_Rdata_ram[59]
  PIN M_Rdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 35.328 0.084 35.352 ;
    END
  END M_Rdata_ram[5]
  PIN M_Rdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.952 0.084 17.976 ;
    END
  END M_Rdata_ram[60]
  PIN M_Rdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.392 0.084 19.416 ;
    END
  END M_Rdata_ram[61]
  PIN M_Rdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.528 0.084 18.552 ;
    END
  END M_Rdata_ram[62]
  PIN M_Rdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.184 41.235 17.208 41.319 ;
    END
  END M_Rdata_ram[63]
  PIN M_Rdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.52 41.235 11.544 41.319 ;
    END
  END M_Rdata_ram[6]
  PIN M_Rdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.328 41.235 11.352 41.319 ;
    END
  END M_Rdata_ram[7]
  PIN M_Rdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.424 0.084 23.448 ;
    END
  END M_Rdata_ram[8]
  PIN M_Rdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.272 0.084 22.296 ;
    END
  END M_Rdata_ram[9]
  PIN Min_Wdata_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 40.32 41.319 40.344 ;
    END
  END Min_Wdata_ram[0]
  PIN Min_Wdata_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.36 41.319 39.384 ;
    END
  END Min_Wdata_ram[10]
  PIN Min_Wdata_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 40.128 41.319 40.152 ;
    END
  END Min_Wdata_ram[11]
  PIN Min_Wdata_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.008 41.235 19.032 41.319 ;
    END
  END Min_Wdata_ram[12]
  PIN Min_Wdata_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.64 0.084 20.664 ;
    END
  END Min_Wdata_ram[13]
  PIN Min_Wdata_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.36 0 39.384 0.084 ;
    END
  END Min_Wdata_ram[14]
  PIN Min_Wdata_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.456 41.319 39.48 ;
    END
  END Min_Wdata_ram[15]
  PIN Min_Wdata_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 40.032 41.319 40.056 ;
    END
  END Min_Wdata_ram[16]
  PIN Min_Wdata_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.84 0 39.864 0.084 ;
    END
  END Min_Wdata_ram[17]
  PIN Min_Wdata_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.176 41.235 10.2 41.319 ;
    END
  END Min_Wdata_ram[18]
  PIN Min_Wdata_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.608 0.084 16.632 ;
    END
  END Min_Wdata_ram[19]
  PIN Min_Wdata_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.792 41.235 33.816 41.319 ;
    END
  END Min_Wdata_ram[1]
  PIN Min_Wdata_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.144 41.235 30.168 41.319 ;
    END
  END Min_Wdata_ram[20]
  PIN Min_Wdata_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.744 0 39.768 0.084 ;
    END
  END Min_Wdata_ram[21]
  PIN Min_Wdata_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.552 0 39.576 0.084 ;
    END
  END Min_Wdata_ram[22]
  PIN Min_Wdata_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.6 41.235 33.624 41.319 ;
    END
  END Min_Wdata_ram[23]
  PIN Min_Wdata_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.92 41.235 1.944 41.319 ;
    END
  END Min_Wdata_ram[24]
  PIN Min_Wdata_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 1.728 0.084 1.752 ;
    END
  END Min_Wdata_ram[25]
  PIN Min_Wdata_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.912 41.235 18.936 41.319 ;
    END
  END Min_Wdata_ram[26]
  PIN Min_Wdata_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.552 41.319 39.576 ;
    END
  END Min_Wdata_ram[27]
  PIN Min_Wdata_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.456 0 39.48 0.084 ;
    END
  END Min_Wdata_ram[28]
  PIN Min_Wdata_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.088 41.235 17.112 41.319 ;
    END
  END Min_Wdata_ram[29]
  PIN Min_Wdata_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.648 0 39.672 0.084 ;
    END
  END Min_Wdata_ram[2]
  PIN Min_Wdata_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.264 41.319 39.288 ;
    END
  END Min_Wdata_ram[30]
  PIN Min_Wdata_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.52 41.319 23.544 ;
    END
  END Min_Wdata_ram[31]
  PIN Min_Wdata_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 31.872 0.084 31.896 ;
    END
  END Min_Wdata_ram[32]
  PIN Min_Wdata_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 31.296 0.084 31.32 ;
    END
  END Min_Wdata_ram[33]
  PIN Min_Wdata_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.432 0.084 30.456 ;
    END
  END Min_Wdata_ram[34]
  PIN Min_Wdata_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.376 0.084 29.4 ;
    END
  END Min_Wdata_ram[35]
  PIN Min_Wdata_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.32 0.084 28.344 ;
    END
  END Min_Wdata_ram[36]
  PIN Min_Wdata_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 27.168 0.084 27.192 ;
    END
  END Min_Wdata_ram[37]
  PIN Min_Wdata_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 26.016 0.084 26.04 ;
    END
  END Min_Wdata_ram[38]
  PIN Min_Wdata_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.864 0.084 24.888 ;
    END
  END Min_Wdata_ram[39]
  PIN Min_Wdata_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.016 41.235 2.04 41.319 ;
    END
  END Min_Wdata_ram[3]
  PIN Min_Wdata_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.808 0.084 23.832 ;
    END
  END Min_Wdata_ram[40]
  PIN Min_Wdata_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.56 0.084 22.584 ;
    END
  END Min_Wdata_ram[41]
  PIN Min_Wdata_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.216 0.084 21.24 ;
    END
  END Min_Wdata_ram[42]
  PIN Min_Wdata_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.256 0.084 20.28 ;
    END
  END Min_Wdata_ram[43]
  PIN Min_Wdata_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.912 0.084 18.936 ;
    END
  END Min_Wdata_ram[44]
  PIN Min_Wdata_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.568 0.084 17.592 ;
    END
  END Min_Wdata_ram[45]
  PIN Min_Wdata_ram[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.128 0.084 16.152 ;
    END
  END Min_Wdata_ram[46]
  PIN Min_Wdata_ram[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.208 0.084 14.232 ;
    END
  END Min_Wdata_ram[47]
  PIN Min_Wdata_ram[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.96 0.084 12.984 ;
    END
  END Min_Wdata_ram[48]
  PIN Min_Wdata_ram[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.944 0.084 10.968 ;
    END
  END Min_Wdata_ram[49]
  PIN Min_Wdata_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.344 41.235 1.368 41.319 ;
    END
  END Min_Wdata_ram[4]
  PIN Min_Wdata_ram[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.08 0.084 10.104 ;
    END
  END Min_Wdata_ram[50]
  PIN Min_Wdata_ram[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.832 0 8.856 0.084 ;
    END
  END Min_Wdata_ram[51]
  PIN Min_Wdata_ram[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.736 0 8.76 0.084 ;
    END
  END Min_Wdata_ram[52]
  PIN Min_Wdata_ram[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.776 0 7.8 0.084 ;
    END
  END Min_Wdata_ram[53]
  PIN Min_Wdata_ram[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.64 0.084 8.664 ;
    END
  END Min_Wdata_ram[54]
  PIN Min_Wdata_ram[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.024 0.084 9.048 ;
    END
  END Min_Wdata_ram[55]
  PIN Min_Wdata_ram[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.312 0.084 9.336 ;
    END
  END Min_Wdata_ram[56]
  PIN Min_Wdata_ram[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.984 0.084 10.008 ;
    END
  END Min_Wdata_ram[57]
  PIN Min_Wdata_ram[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.328 0.084 11.352 ;
    END
  END Min_Wdata_ram[58]
  PIN Min_Wdata_ram[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.384 0.084 12.408 ;
    END
  END Min_Wdata_ram[59]
  PIN Min_Wdata_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.096 0 24.12 0.084 ;
    END
  END Min_Wdata_ram[5]
  PIN Min_Wdata_ram[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.768 0.084 12.792 ;
    END
  END Min_Wdata_ram[60]
  PIN Min_Wdata_ram[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.824 0.084 13.848 ;
    END
  END Min_Wdata_ram[61]
  PIN Min_Wdata_ram[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.88 0.084 14.904 ;
    END
  END Min_Wdata_ram[62]
  PIN Min_Wdata_ram[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.624 0.084 30.648 ;
    END
  END Min_Wdata_ram[63]
  PIN Min_Wdata_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.992 41.235 17.016 41.319 ;
    END
  END Min_Wdata_ram[6]
  PIN Min_Wdata_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.072 0 39.096 0.084 ;
    END
  END Min_Wdata_ram[7]
  PIN Min_Wdata_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 29.184 41.319 29.208 ;
    END
  END Min_Wdata_ram[8]
  PIN Min_Wdata_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 18.624 41.319 18.648 ;
    END
  END Min_Wdata_ram[9]
  PIN Min_addr_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.592 41.235 14.616 41.319 ;
    END
  END Min_addr_ram[0]
  PIN Min_addr_ram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.096 41.235 12.12 41.319 ;
    END
  END Min_addr_ram[10]
  PIN Min_addr_ram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.128 41.235 16.152 41.319 ;
    END
  END Min_addr_ram[11]
  PIN Min_addr_ram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.68 0.084 19.704 ;
    END
  END Min_addr_ram[12]
  PIN Min_addr_ram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.856 0.084 17.88 ;
    END
  END Min_addr_ram[13]
  PIN Min_addr_ram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.32 0.084 16.344 ;
    END
  END Min_addr_ram[14]
  PIN Min_addr_ram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.456 0.084 15.48 ;
    END
  END Min_addr_ram[15]
  PIN Min_addr_ram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.84 0.084 15.864 ;
    END
  END Min_addr_ram[16]
  PIN Min_addr_ram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.384 0 12.408 0.084 ;
    END
  END Min_addr_ram[17]
  PIN Min_addr_ram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.032 0 16.056 0.084 ;
    END
  END Min_addr_ram[18]
  PIN Min_addr_ram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.88 0 14.904 0.084 ;
    END
  END Min_addr_ram[19]
  PIN Min_addr_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.688 41.235 14.712 41.319 ;
    END
  END Min_addr_ram[1]
  PIN Min_addr_ram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.936 0 15.96 0.084 ;
    END
  END Min_addr_ram[20]
  PIN Min_addr_ram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.248 0 13.272 0.084 ;
    END
  END Min_addr_ram[21]
  PIN Min_addr_ram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.744 41.235 15.768 41.319 ;
    END
  END Min_addr_ram[22]
  PIN Min_addr_ram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.136 41.235 23.16 41.319 ;
    END
  END Min_addr_ram[23]
  PIN Min_addr_ram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.216 41.235 21.24 41.319 ;
    END
  END Min_addr_ram[24]
  PIN Min_addr_ram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.08 41.235 22.104 41.319 ;
    END
  END Min_addr_ram[25]
  PIN Min_addr_ram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 41.235 21.72 41.319 ;
    END
  END Min_addr_ram[26]
  PIN Min_addr_ram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.896 41.319 28.92 ;
    END
  END Min_addr_ram[27]
  PIN Min_addr_ram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.128 41.319 28.152 ;
    END
  END Min_addr_ram[28]
  PIN Min_addr_ram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 26.016 41.319 26.04 ;
    END
  END Min_addr_ram[29]
  PIN Min_addr_ram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.168 41.235 15.192 41.319 ;
    END
  END Min_addr_ram[2]
  PIN Min_addr_ram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.632 41.319 25.656 ;
    END
  END Min_addr_ram[30]
  PIN Min_addr_ram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 24.384 41.319 24.408 ;
    END
  END Min_addr_ram[31]
  PIN Min_addr_ram[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.232 41.319 23.256 ;
    END
  END Min_addr_ram[32]
  PIN Min_addr_ram[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 21.984 41.319 22.008 ;
    END
  END Min_addr_ram[33]
  PIN Min_addr_ram[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 20.736 41.319 20.76 ;
    END
  END Min_addr_ram[34]
  PIN Min_addr_ram[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.312 0 21.336 0.084 ;
    END
  END Min_addr_ram[35]
  PIN Min_addr_ram[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 0 21.72 0.084 ;
    END
  END Min_addr_ram[36]
  PIN Min_addr_ram[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.792 0 21.816 0.084 ;
    END
  END Min_addr_ram[37]
  PIN Min_addr_ram[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.272 0 22.296 0.084 ;
    END
  END Min_addr_ram[38]
  PIN Min_addr_ram[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.56 0 22.584 0.084 ;
    END
  END Min_addr_ram[39]
  PIN Min_addr_ram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.288 41.235 12.312 41.319 ;
    END
  END Min_addr_ram[3]
  PIN Min_addr_ram[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 0 22.008 0.084 ;
    END
  END Min_addr_ram[40]
  PIN Min_addr_ram[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.752 0 22.776 0.084 ;
    END
  END Min_addr_ram[41]
  PIN Min_addr_ram[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.368 0 22.392 0.084 ;
    END
  END Min_addr_ram[42]
  PIN Min_addr_ram[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.544 0 20.568 0.084 ;
    END
  END Min_addr_ram[43]
  PIN Min_addr_ram[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.848 0 22.872 0.084 ;
    END
  END Min_addr_ram[44]
  PIN Min_addr_ram[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.344 41.319 25.368 ;
    END
  END Min_addr_ram[45]
  PIN Min_addr_ram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.976 41.235 15 41.319 ;
    END
  END Min_addr_ram[4]
  PIN Min_addr_ram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.072 41.235 15.096 41.319 ;
    END
  END Min_addr_ram[5]
  PIN Min_addr_ram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.648 41.235 15.672 41.319 ;
    END
  END Min_addr_ram[6]
  PIN Min_addr_ram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.84 41.235 15.864 41.319 ;
    END
  END Min_addr_ram[7]
  PIN Min_addr_ram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.32 41.235 16.344 41.319 ;
    END
  END Min_addr_ram[8]
  PIN Min_addr_ram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.192 41.235 12.216 41.319 ;
    END
  END Min_addr_ram[9]
  PIN Min_data_ram_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.144 41.235 18.168 41.319 ;
    END
  END Min_data_ram_size[0]
  PIN Min_data_ram_size[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.328 0 23.352 0.084 ;
    END
  END Min_data_ram_size[10]
  PIN Min_data_ram_size[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.544 41.235 20.568 41.319 ;
    END
  END Min_data_ram_size[11]
  PIN Min_data_ram_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.856 41.235 17.88 41.319 ;
    END
  END Min_data_ram_size[1]
  PIN Min_data_ram_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.048 41.235 18.072 41.319 ;
    END
  END Min_data_ram_size[2]
  PIN Min_data_ram_size[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.512 41.235 16.536 41.319 ;
    END
  END Min_data_ram_size[3]
  PIN Min_data_ram_size[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  17.952 41.235 17.976 41.319 ;
    END
  END Min_data_ram_size[4]
  PIN Min_data_ram_size[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.24 41.235 18.264 41.319 ;
    END
  END Min_data_ram_size[5]
  PIN Min_data_ram_size[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.712 0 23.736 0.084 ;
    END
  END Min_data_ram_size[6]
  PIN Min_data_ram_size[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.136 0 23.16 0.084 ;
    END
  END Min_data_ram_size[7]
  PIN Min_data_ram_size[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.232 0 23.256 0.084 ;
    END
  END Min_data_ram_size[8]
  PIN Min_data_ram_size[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.448 41.235 20.472 41.319 ;
    END
  END Min_data_ram_size[9]
  PIN Min_oe_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.032 41.235 16.056 41.319 ;
    END
  END Min_oe_ram[0]
  PIN Min_oe_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.408 41.235 21.432 41.319 ;
    END
  END Min_oe_ram[1]
  PIN Min_we_ram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 34.848 0.084 34.872 ;
    END
  END Min_we_ram[0]
  PIN Min_we_ram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.8 0 16.824 0.084 ;
    END
  END Min_we_ram[1]
  PIN Mout_Wdata_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.648 41.319 39.672 ;
    END
  END Mout_Wdata_ram[0]
  PIN Mout_Wdata_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.072 41.319 39.096 ;
    END
  END Mout_Wdata_ram[10]
  PIN Mout_Wdata_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.84 41.319 39.864 ;
    END
  END Mout_Wdata_ram[11]
  PIN Mout_Wdata_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.2 41.235 19.224 41.319 ;
    END
  END Mout_Wdata_ram[12]
  PIN Mout_Wdata_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.544 0.084 20.568 ;
    END
  END Mout_Wdata_ram[13]
  PIN Mout_Wdata_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.264 0 39.288 0.084 ;
    END
  END Mout_Wdata_ram[14]
  PIN Mout_Wdata_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.744 41.319 39.768 ;
    END
  END Mout_Wdata_ram[15]
  PIN Mout_Wdata_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 40.224 41.319 40.248 ;
    END
  END Mout_Wdata_ram[16]
  PIN Mout_Wdata_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.32 0 40.344 0.084 ;
    END
  END Mout_Wdata_ram[17]
  PIN Mout_Wdata_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.368 41.235 10.392 41.319 ;
    END
  END Mout_Wdata_ram[18]
  PIN Mout_Wdata_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.704 0.084 16.728 ;
    END
  END Mout_Wdata_ram[19]
  PIN Mout_Wdata_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.984 41.235 34.008 41.319 ;
    END
  END Mout_Wdata_ram[1]
  PIN Mout_Wdata_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.336 41.235 30.36 41.319 ;
    END
  END Mout_Wdata_ram[20]
  PIN Mout_Wdata_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.224 0 40.248 0.084 ;
    END
  END Mout_Wdata_ram[21]
  PIN Mout_Wdata_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.032 0 40.056 0.084 ;
    END
  END Mout_Wdata_ram[22]
  PIN Mout_Wdata_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.696 41.235 33.72 41.319 ;
    END
  END Mout_Wdata_ram[23]
  PIN Mout_Wdata_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.112 41.235 2.136 41.319 ;
    END
  END Mout_Wdata_ram[24]
  PIN Mout_Wdata_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 1.632 0.084 1.656 ;
    END
  END Mout_Wdata_ram[25]
  PIN Mout_Wdata_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.104 41.235 19.128 41.319 ;
    END
  END Mout_Wdata_ram[26]
  PIN Mout_Wdata_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.168 41.319 39.192 ;
    END
  END Mout_Wdata_ram[27]
  PIN Mout_Wdata_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.936 0 39.96 0.084 ;
    END
  END Mout_Wdata_ram[28]
  PIN Mout_Wdata_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.8 41.235 16.824 41.319 ;
    END
  END Mout_Wdata_ram[29]
  PIN Mout_Wdata_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  40.128 0 40.152 0.084 ;
    END
  END Mout_Wdata_ram[2]
  PIN Mout_Wdata_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 39.936 41.319 39.96 ;
    END
  END Mout_Wdata_ram[30]
  PIN Mout_Wdata_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.616 41.319 23.64 ;
    END
  END Mout_Wdata_ram[31]
  PIN Mout_Wdata_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 31.776 0.084 31.8 ;
    END
  END Mout_Wdata_ram[32]
  PIN Mout_Wdata_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 31.392 0.084 31.416 ;
    END
  END Mout_Wdata_ram[33]
  PIN Mout_Wdata_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.336 0.084 30.36 ;
    END
  END Mout_Wdata_ram[34]
  PIN Mout_Wdata_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.28 0.084 29.304 ;
    END
  END Mout_Wdata_ram[35]
  PIN Mout_Wdata_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.224 0.084 28.248 ;
    END
  END Mout_Wdata_ram[36]
  PIN Mout_Wdata_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 27.072 0.084 27.096 ;
    END
  END Mout_Wdata_ram[37]
  PIN Mout_Wdata_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.92 0.084 25.944 ;
    END
  END Mout_Wdata_ram[38]
  PIN Mout_Wdata_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.768 0.084 24.792 ;
    END
  END Mout_Wdata_ram[39]
  PIN Mout_Wdata_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.208 41.235 2.232 41.319 ;
    END
  END Mout_Wdata_ram[3]
  PIN Mout_Wdata_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.712 0.084 23.736 ;
    END
  END Mout_Wdata_ram[40]
  PIN Mout_Wdata_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 22.464 0.084 22.488 ;
    END
  END Mout_Wdata_ram[41]
  PIN Mout_Wdata_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.12 0.084 21.144 ;
    END
  END Mout_Wdata_ram[42]
  PIN Mout_Wdata_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.16 0.084 20.184 ;
    END
  END Mout_Wdata_ram[43]
  PIN Mout_Wdata_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.816 0.084 18.84 ;
    END
  END Mout_Wdata_ram[44]
  PIN Mout_Wdata_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.472 0.084 17.496 ;
    END
  END Mout_Wdata_ram[45]
  PIN Mout_Wdata_ram[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.032 0.084 16.056 ;
    END
  END Mout_Wdata_ram[46]
  PIN Mout_Wdata_ram[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.304 0.084 14.328 ;
    END
  END Mout_Wdata_ram[47]
  PIN Mout_Wdata_ram[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.864 0.084 12.888 ;
    END
  END Mout_Wdata_ram[48]
  PIN Mout_Wdata_ram[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.848 0.084 10.872 ;
    END
  END Mout_Wdata_ram[49]
  PIN Mout_Wdata_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.536 41.235 1.56 41.319 ;
    END
  END Mout_Wdata_ram[4]
  PIN Mout_Wdata_ram[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.792 0.084 9.816 ;
    END
  END Mout_Wdata_ram[50]
  PIN Mout_Wdata_ram[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.12 0 9.144 0.084 ;
    END
  END Mout_Wdata_ram[51]
  PIN Mout_Wdata_ram[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.024 0 9.048 0.084 ;
    END
  END Mout_Wdata_ram[52]
  PIN Mout_Wdata_ram[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.064 0 8.088 0.084 ;
    END
  END Mout_Wdata_ram[53]
  PIN Mout_Wdata_ram[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.544 0.084 8.568 ;
    END
  END Mout_Wdata_ram[54]
  PIN Mout_Wdata_ram[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.928 0.084 8.952 ;
    END
  END Mout_Wdata_ram[55]
  PIN Mout_Wdata_ram[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.216 0.084 9.24 ;
    END
  END Mout_Wdata_ram[56]
  PIN Mout_Wdata_ram[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.888 0.084 9.912 ;
    END
  END Mout_Wdata_ram[57]
  PIN Mout_Wdata_ram[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.232 0.084 11.256 ;
    END
  END Mout_Wdata_ram[58]
  PIN Mout_Wdata_ram[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.288 0.084 12.312 ;
    END
  END Mout_Wdata_ram[59]
  PIN Mout_Wdata_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.808 0 23.832 0.084 ;
    END
  END Mout_Wdata_ram[5]
  PIN Mout_Wdata_ram[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.672 0.084 12.696 ;
    END
  END Mout_Wdata_ram[60]
  PIN Mout_Wdata_ram[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.728 0.084 13.752 ;
    END
  END Mout_Wdata_ram[61]
  PIN Mout_Wdata_ram[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.784 0.084 14.808 ;
    END
  END Mout_Wdata_ram[62]
  PIN Mout_Wdata_ram[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.528 0.084 30.552 ;
    END
  END Mout_Wdata_ram[63]
  PIN Mout_Wdata_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.896 41.235 16.92 41.319 ;
    END
  END Mout_Wdata_ram[6]
  PIN Mout_Wdata_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  39.168 0 39.192 0.084 ;
    END
  END Mout_Wdata_ram[7]
  PIN Mout_Wdata_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 29.088 41.319 29.112 ;
    END
  END Mout_Wdata_ram[8]
  PIN Mout_Wdata_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 18.72 41.319 18.744 ;
    END
  END Mout_Wdata_ram[9]
  PIN Mout_addr_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.784 41.235 14.808 41.319 ;
    END
  END Mout_addr_ram[0]
  PIN Mout_addr_ram[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.904 41.235 11.928 41.319 ;
    END
  END Mout_addr_ram[10]
  PIN Mout_addr_ram[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.416 41.235 16.44 41.319 ;
    END
  END Mout_addr_ram[11]
  PIN Mout_addr_ram[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.584 0.084 19.608 ;
    END
  END Mout_addr_ram[12]
  PIN Mout_addr_ram[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.76 0.084 17.784 ;
    END
  END Mout_addr_ram[13]
  PIN Mout_addr_ram[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.224 0.084 16.248 ;
    END
  END Mout_addr_ram[14]
  PIN Mout_addr_ram[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.36 0.084 15.384 ;
    END
  END Mout_addr_ram[15]
  PIN Mout_addr_ram[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.936 0.084 15.96 ;
    END
  END Mout_addr_ram[16]
  PIN Mout_addr_ram[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.672 0 12.696 0.084 ;
    END
  END Mout_addr_ram[17]
  PIN Mout_addr_ram[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.32 0 16.344 0.084 ;
    END
  END Mout_addr_ram[18]
  PIN Mout_addr_ram[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.168 0 15.192 0.084 ;
    END
  END Mout_addr_ram[19]
  PIN Mout_addr_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  14.88 41.235 14.904 41.319 ;
    END
  END Mout_addr_ram[1]
  PIN Mout_addr_ram[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.224 0 16.248 0.084 ;
    END
  END Mout_addr_ram[20]
  PIN Mout_addr_ram[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.536 0 13.56 0.084 ;
    END
  END Mout_addr_ram[21]
  PIN Mout_addr_ram[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  13.632 0 13.656 0.084 ;
    END
  END Mout_addr_ram[22]
  PIN Mout_addr_ram[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.424 41.235 23.448 41.319 ;
    END
  END Mout_addr_ram[23]
  PIN Mout_addr_ram[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.6 41.235 21.624 41.319 ;
    END
  END Mout_addr_ram[24]
  PIN Mout_addr_ram[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.368 41.235 22.392 41.319 ;
    END
  END Mout_addr_ram[25]
  PIN Mout_addr_ram[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 41.235 22.008 41.319 ;
    END
  END Mout_addr_ram[26]
  PIN Mout_addr_ram[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.992 41.319 29.016 ;
    END
  END Mout_addr_ram[27]
  PIN Mout_addr_ram[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.032 41.319 28.056 ;
    END
  END Mout_addr_ram[28]
  PIN Mout_addr_ram[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.92 41.319 25.944 ;
    END
  END Mout_addr_ram[29]
  PIN Mout_addr_ram[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.456 41.235 15.48 41.319 ;
    END
  END Mout_addr_ram[2]
  PIN Mout_addr_ram[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.536 41.319 25.56 ;
    END
  END Mout_addr_ram[30]
  PIN Mout_addr_ram[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 24.48 41.319 24.504 ;
    END
  END Mout_addr_ram[31]
  PIN Mout_addr_ram[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.328 41.319 23.352 ;
    END
  END Mout_addr_ram[32]
  PIN Mout_addr_ram[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 22.08 41.319 22.104 ;
    END
  END Mout_addr_ram[33]
  PIN Mout_addr_ram[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 20.832 41.319 20.856 ;
    END
  END Mout_addr_ram[34]
  PIN Mout_addr_ram[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.504 0 21.528 0.084 ;
    END
  END Mout_addr_ram[35]
  PIN Mout_addr_ram[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.888 0 21.912 0.084 ;
    END
  END Mout_addr_ram[36]
  PIN Mout_addr_ram[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.08 0 22.104 0.084 ;
    END
  END Mout_addr_ram[37]
  PIN Mout_addr_ram[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.464 0 22.488 0.084 ;
    END
  END Mout_addr_ram[38]
  PIN Mout_addr_ram[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.04 0 23.064 0.084 ;
    END
  END Mout_addr_ram[39]
  PIN Mout_addr_ram[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.576 41.235 12.6 41.319 ;
    END
  END Mout_addr_ram[3]
  PIN Mout_addr_ram[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.176 0 22.2 0.084 ;
    END
  END Mout_addr_ram[40]
  PIN Mout_addr_ram[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.944 0 22.968 0.084 ;
    END
  END Mout_addr_ram[41]
  PIN Mout_addr_ram[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.656 0 22.68 0.084 ;
    END
  END Mout_addr_ram[42]
  PIN Mout_addr_ram[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.832 0 20.856 0.084 ;
    END
  END Mout_addr_ram[43]
  PIN Mout_addr_ram[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24 0 24.024 0.084 ;
    END
  END Mout_addr_ram[44]
  PIN Mout_addr_ram[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.248 41.319 25.272 ;
    END
  END Mout_addr_ram[45]
  PIN Mout_addr_ram[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.264 41.235 15.288 41.319 ;
    END
  END Mout_addr_ram[4]
  PIN Mout_addr_ram[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.36 41.235 15.384 41.319 ;
    END
  END Mout_addr_ram[5]
  PIN Mout_addr_ram[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.552 41.235 15.576 41.319 ;
    END
  END Mout_addr_ram[6]
  PIN Mout_addr_ram[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.936 41.235 15.96 41.319 ;
    END
  END Mout_addr_ram[7]
  PIN Mout_addr_ram[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.608 41.235 16.632 41.319 ;
    END
  END Mout_addr_ram[8]
  PIN Mout_addr_ram[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  12.48 41.235 12.504 41.319 ;
    END
  END Mout_addr_ram[9]
  PIN Mout_data_ram_size[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.72 41.235 18.744 41.319 ;
    END
  END Mout_data_ram_size[0]
  PIN Mout_data_ram_size[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.52 0 23.544 0.084 ;
    END
  END Mout_data_ram_size[10]
  PIN Mout_data_ram_size[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.64 41.235 20.664 41.319 ;
    END
  END Mout_data_ram_size[11]
  PIN Mout_data_ram_size[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.336 41.235 18.36 41.319 ;
    END
  END Mout_data_ram_size[1]
  PIN Mout_data_ram_size[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.432 41.235 18.456 41.319 ;
    END
  END Mout_data_ram_size[2]
  PIN Mout_data_ram_size[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.704 41.235 16.728 41.319 ;
    END
  END Mout_data_ram_size[3]
  PIN Mout_data_ram_size[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.528 41.235 18.552 41.319 ;
    END
  END Mout_data_ram_size[4]
  PIN Mout_data_ram_size[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  18.624 41.235 18.648 41.319 ;
    END
  END Mout_data_ram_size[5]
  PIN Mout_data_ram_size[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.904 0 23.928 0.084 ;
    END
  END Mout_data_ram_size[6]
  PIN Mout_data_ram_size[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.616 0 23.64 0.084 ;
    END
  END Mout_data_ram_size[7]
  PIN Mout_data_ram_size[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.424 0 23.448 0.084 ;
    END
  END Mout_data_ram_size[8]
  PIN Mout_data_ram_size[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.736 41.235 20.76 41.319 ;
    END
  END Mout_data_ram_size[9]
  PIN Mout_oe_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.224 41.235 16.248 41.319 ;
    END
  END Mout_oe_ram[0]
  PIN Mout_oe_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.12 41.235 21.144 41.319 ;
    END
  END Mout_oe_ram[1]
  PIN Mout_we_ram[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 34.944 0.084 34.968 ;
    END
  END Mout_we_ram[0]
  PIN Mout_we_ram[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  16.992 0 17.016 0.084 ;
    END
  END Mout_we_ram[1]
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  36.288 41.235 36.312 41.319 ;
    END
  END clock
  PIN done_port
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.36 41.235 27.384 41.319 ;
    END
  END done_port
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.312 41.235 21.336 41.319 ;
    END
  END reset
  PIN start_port
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  27.168 41.235 27.192 41.319 ;
    END
  END start_port
  PIN vargs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  29.376 41.235 29.4 41.319 ;
    END
  END vargs[0]
  PIN vargs[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 20.64 41.319 20.664 ;
    END
  END vargs[10]
  PIN vargs[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 19.872 41.319 19.896 ;
    END
  END vargs[11]
  PIN vargs[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 14.88 41.319 14.904 ;
    END
  END vargs[12]
  PIN vargs[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 14.4 41.319 14.424 ;
    END
  END vargs[13]
  PIN vargs[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 14.016 41.319 14.04 ;
    END
  END vargs[14]
  PIN vargs[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 14.112 41.319 14.136 ;
    END
  END vargs[15]
  PIN vargs[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 12.768 41.319 12.792 ;
    END
  END vargs[16]
  PIN vargs[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 11.136 41.319 11.16 ;
    END
  END vargs[17]
  PIN vargs[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 10.848 41.319 10.872 ;
    END
  END vargs[18]
  PIN vargs[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 10.944 41.319 10.968 ;
    END
  END vargs[19]
  PIN vargs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.976 41.235 27 41.319 ;
    END
  END vargs[1]
  PIN vargs[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.992 0 29.016 0.084 ;
    END
  END vargs[20]
  PIN vargs[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  28.32 0 28.344 0.084 ;
    END
  END vargs[21]
  PIN vargs[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.048 0 30.072 0.084 ;
    END
  END vargs[22]
  PIN vargs[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.432 0 30.456 0.084 ;
    END
  END vargs[23]
  PIN vargs[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.528 0 30.552 0.084 ;
    END
  END vargs[24]
  PIN vargs[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  30.624 0 30.648 0.084 ;
    END
  END vargs[25]
  PIN vargs[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.296 0 31.32 0.084 ;
    END
  END vargs[26]
  PIN vargs[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.584 0 31.608 0.084 ;
    END
  END vargs[27]
  PIN vargs[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  31.872 0 31.896 0.084 ;
    END
  END vargs[28]
  PIN vargs[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.544 0 32.568 0.084 ;
    END
  END vargs[29]
  PIN vargs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.224 41.319 28.248 ;
    END
  END vargs[2]
  PIN vargs[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  32.832 0 32.856 0.084 ;
    END
  END vargs[30]
  PIN vargs[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  33.504 0 33.528 0.084 ;
    END
  END vargs[31]
  PIN vargs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 28.32 41.319 28.344 ;
    END
  END vargs[3]
  PIN vargs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 27.744 41.319 27.768 ;
    END
  END vargs[4]
  PIN vargs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 25.728 41.319 25.752 ;
    END
  END vargs[5]
  PIN vargs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 24.096 41.319 24.12 ;
    END
  END vargs[6]
  PIN vargs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.712 41.319 23.736 ;
    END
  END vargs[7]
  PIN vargs[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.808 41.319 23.832 ;
    END
  END vargs[8]
  PIN vargs[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  41.235 23.136 41.319 23.16 ;
    END
  END vargs[9]
  OBS
    LAYER M1 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M2 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M3 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M4 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M5 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M6 ;
     RECT  0 0 41.319 41.319 ;
    LAYER M7 ;
     RECT  0 0 41.319 41.319 ;
  END
END run_benchmark
END LIBRARY
