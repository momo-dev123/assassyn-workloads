VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA pe_5_2_via1_2_10692_18_1_297_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 297 ;
END pe_5_2_via1_2_10692_18_1_297_36_36

VIA pe_5_2_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END pe_5_2_VIA23_1_3_36_36

VIA pe_5_2_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END pe_5_2_VIA34_1_2_58_52

VIA pe_5_2_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END pe_5_2_VIA45_1_2_58_58

VIA pe_5_2_via5_6_120_288_1_2_58_322
  VIARULE M6_M5widePWR1p152 ;
  CUTSIZE 0.024 0.288 ;
  LAYERS M5 V5 M6 ;
  CUTSPACING 0.034 0.034 ;
  ENCLOSURE 0.019 0 0 0 ;
  ROWCOL 1 2 ;
END pe_5_2_via5_6_120_288_1_2_58_322

MACRO pe_5_2
  FOREIGN pe_5_2 0 0 ;
  CLASS BLOCK ;
  SIZE 12.737 BY 12.737 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.458 7.833 7.482 8.121 ;
        RECT  1.458 1.833 7.482 2.121 ;
      LAYER M5 ;
        RECT  7.362 1.327 7.482 11.633 ;
        RECT  1.458 1.327 1.578 11.633 ;
      LAYER M2 ;
        RECT  1.026 11.601 11.718 11.619 ;
        RECT  1.026 11.061 11.718 11.079 ;
        RECT  1.026 10.521 11.718 10.539 ;
        RECT  1.026 9.981 11.718 9.999 ;
        RECT  1.026 9.441 11.718 9.459 ;
        RECT  1.026 8.901 11.718 8.919 ;
        RECT  1.026 8.361 11.718 8.379 ;
        RECT  1.026 7.821 11.718 7.839 ;
        RECT  1.026 7.281 11.718 7.299 ;
        RECT  1.026 6.741 11.718 6.759 ;
        RECT  1.026 6.201 11.718 6.219 ;
        RECT  1.026 5.661 11.718 5.679 ;
        RECT  1.026 5.121 11.718 5.139 ;
        RECT  1.026 4.581 11.718 4.599 ;
        RECT  1.026 4.041 11.718 4.059 ;
        RECT  1.026 3.501 11.718 3.519 ;
        RECT  1.026 2.961 11.718 2.979 ;
        RECT  1.026 2.421 11.718 2.439 ;
        RECT  1.026 1.881 11.718 1.899 ;
        RECT  1.026 1.341 11.718 1.359 ;
      LAYER M1 ;
        RECT  1.026 11.601 11.718 11.619 ;
        RECT  1.026 11.061 11.718 11.079 ;
        RECT  1.026 10.521 11.718 10.539 ;
        RECT  1.026 9.981 11.718 9.999 ;
        RECT  1.026 9.441 11.718 9.459 ;
        RECT  1.026 8.901 11.718 8.919 ;
        RECT  1.026 8.361 11.718 8.379 ;
        RECT  1.026 7.821 11.718 7.839 ;
        RECT  1.026 7.281 11.718 7.299 ;
        RECT  1.026 6.741 11.718 6.759 ;
        RECT  1.026 6.201 11.718 6.219 ;
        RECT  1.026 5.661 11.718 5.679 ;
        RECT  1.026 5.121 11.718 5.139 ;
        RECT  1.026 4.581 11.718 4.599 ;
        RECT  1.026 4.041 11.718 4.059 ;
        RECT  1.026 3.501 11.718 3.519 ;
        RECT  1.026 2.961 11.718 2.979 ;
        RECT  1.026 2.421 11.718 2.439 ;
        RECT  1.026 1.881 11.718 1.899 ;
        RECT  1.026 1.341 11.718 1.359 ;
      VIA 7.422 7.977 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 1.977 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 7.977 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 1.518 1.977 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 7.422 11.61 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.593 7.467 11.627 ;
      VIA 7.422 11.61 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 11.61 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 11.07 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 11.053 7.467 11.087 ;
      VIA 7.422 11.07 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 11.07 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 10.53 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 10.513 7.467 10.547 ;
      VIA 7.422 10.53 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 10.53 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 9.99 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.973 7.467 10.007 ;
      VIA 7.422 9.99 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 9.99 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 9.45 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 9.433 7.467 9.467 ;
      VIA 7.422 9.45 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 9.45 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 8.91 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.893 7.467 8.927 ;
      VIA 7.422 8.91 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 8.91 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 8.37 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 8.353 7.467 8.387 ;
      VIA 7.422 8.37 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 8.37 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 7.83 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.813 7.467 7.847 ;
      VIA 7.422 7.83 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 7.83 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 7.29 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 7.273 7.467 7.307 ;
      VIA 7.422 7.29 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 7.29 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 6.75 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.733 7.467 6.767 ;
      VIA 7.422 6.75 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 6.75 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 6.21 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 6.193 7.467 6.227 ;
      VIA 7.422 6.21 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 6.21 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 5.67 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.653 7.467 5.687 ;
      VIA 7.422 5.67 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 5.67 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 5.13 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 5.113 7.467 5.147 ;
      VIA 7.422 5.13 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 5.13 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 4.59 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.573 7.467 4.607 ;
      VIA 7.422 4.59 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 4.59 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 4.05 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 4.033 7.467 4.067 ;
      VIA 7.422 4.05 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 4.05 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 3.51 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 3.493 7.467 3.527 ;
      VIA 7.422 3.51 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 3.51 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 2.97 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.953 7.467 2.987 ;
      VIA 7.422 2.97 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 2.97 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 2.43 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 2.413 7.467 2.447 ;
      VIA 7.422 2.43 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 2.43 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 1.89 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.873 7.467 1.907 ;
      VIA 7.422 1.89 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 1.89 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.422 1.35 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.377 1.333 7.467 1.367 ;
      VIA 7.422 1.35 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.422 1.35 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 11.61 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.593 1.563 11.627 ;
      VIA 1.518 11.61 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 11.61 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 11.07 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 11.053 1.563 11.087 ;
      VIA 1.518 11.07 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 11.07 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 10.53 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 10.513 1.563 10.547 ;
      VIA 1.518 10.53 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 10.53 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 9.99 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.973 1.563 10.007 ;
      VIA 1.518 9.99 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 9.99 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 9.45 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 9.433 1.563 9.467 ;
      VIA 1.518 9.45 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 9.45 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 8.91 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.893 1.563 8.927 ;
      VIA 1.518 8.91 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 8.91 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 8.37 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 8.353 1.563 8.387 ;
      VIA 1.518 8.37 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 8.37 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 7.83 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.813 1.563 7.847 ;
      VIA 1.518 7.83 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 7.83 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 7.29 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 7.273 1.563 7.307 ;
      VIA 1.518 7.29 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 7.29 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 6.75 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.733 1.563 6.767 ;
      VIA 1.518 6.75 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 6.75 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 6.21 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 6.193 1.563 6.227 ;
      VIA 1.518 6.21 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 6.21 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 5.67 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.653 1.563 5.687 ;
      VIA 1.518 5.67 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 5.67 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 5.13 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 5.113 1.563 5.147 ;
      VIA 1.518 5.13 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 5.13 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 4.59 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.573 1.563 4.607 ;
      VIA 1.518 4.59 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 4.59 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 4.05 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 4.033 1.563 4.067 ;
      VIA 1.518 4.05 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 4.05 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 3.51 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 3.493 1.563 3.527 ;
      VIA 1.518 3.51 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 3.51 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 2.97 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.953 1.563 2.987 ;
      VIA 1.518 2.97 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 2.97 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 2.43 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 2.413 1.563 2.447 ;
      VIA 1.518 2.43 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 2.43 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 1.89 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.873 1.563 1.907 ;
      VIA 1.518 1.89 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 1.89 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.518 1.35 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.473 1.333 1.563 1.367 ;
      VIA 1.518 1.35 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.518 1.35 pe_5_2_VIA23_1_3_36_36 ;
      VIA 6.372 11.61 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 11.07 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 10.53 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 9.99 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 9.45 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 8.91 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 8.37 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 7.83 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 7.29 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 6.75 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 6.21 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 5.67 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 5.13 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 4.59 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 4.05 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 3.51 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 2.97 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 2.43 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 1.89 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 1.35 pe_5_2_via1_2_10692_18_1_297_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M6 ;
        RECT  1.266 7.449 7.29 7.737 ;
        RECT  1.266 1.449 7.29 1.737 ;
      LAYER M5 ;
        RECT  7.17 1.057 7.29 11.363 ;
        RECT  1.266 1.057 1.386 11.363 ;
      LAYER M2 ;
        RECT  1.026 11.331 11.718 11.349 ;
        RECT  1.026 10.791 11.718 10.809 ;
        RECT  1.026 10.251 11.718 10.269 ;
        RECT  1.026 9.711 11.718 9.729 ;
        RECT  1.026 9.171 11.718 9.189 ;
        RECT  1.026 8.631 11.718 8.649 ;
        RECT  1.026 8.091 11.718 8.109 ;
        RECT  1.026 7.551 11.718 7.569 ;
        RECT  1.026 7.011 11.718 7.029 ;
        RECT  1.026 6.471 11.718 6.489 ;
        RECT  1.026 5.931 11.718 5.949 ;
        RECT  1.026 5.391 11.718 5.409 ;
        RECT  1.026 4.851 11.718 4.869 ;
        RECT  1.026 4.311 11.718 4.329 ;
        RECT  1.026 3.771 11.718 3.789 ;
        RECT  1.026 3.231 11.718 3.249 ;
        RECT  1.026 2.691 11.718 2.709 ;
        RECT  1.026 2.151 11.718 2.169 ;
        RECT  1.026 1.611 11.718 1.629 ;
        RECT  1.026 1.071 11.718 1.089 ;
      LAYER M1 ;
        RECT  1.026 11.331 11.718 11.349 ;
        RECT  1.026 10.791 11.718 10.809 ;
        RECT  1.026 10.251 11.718 10.269 ;
        RECT  1.026 9.711 11.718 9.729 ;
        RECT  1.026 9.171 11.718 9.189 ;
        RECT  1.026 8.631 11.718 8.649 ;
        RECT  1.026 8.091 11.718 8.109 ;
        RECT  1.026 7.551 11.718 7.569 ;
        RECT  1.026 7.011 11.718 7.029 ;
        RECT  1.026 6.471 11.718 6.489 ;
        RECT  1.026 5.931 11.718 5.949 ;
        RECT  1.026 5.391 11.718 5.409 ;
        RECT  1.026 4.851 11.718 4.869 ;
        RECT  1.026 4.311 11.718 4.329 ;
        RECT  1.026 3.771 11.718 3.789 ;
        RECT  1.026 3.231 11.718 3.249 ;
        RECT  1.026 2.691 11.718 2.709 ;
        RECT  1.026 2.151 11.718 2.169 ;
        RECT  1.026 1.611 11.718 1.629 ;
        RECT  1.026 1.071 11.718 1.089 ;
      VIA 7.23 7.593 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 1.593 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 7.593 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 1.326 1.593 pe_5_2_via5_6_120_288_1_2_58_322 ;
      VIA 7.23 11.34 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 11.323 7.275 11.357 ;
      VIA 7.23 11.34 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 11.34 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 10.8 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.783 7.275 10.817 ;
      VIA 7.23 10.8 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 10.8 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 10.26 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 10.243 7.275 10.277 ;
      VIA 7.23 10.26 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 10.26 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 9.72 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.703 7.275 9.737 ;
      VIA 7.23 9.72 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 9.72 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 9.18 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 9.163 7.275 9.197 ;
      VIA 7.23 9.18 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 9.18 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 8.64 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.623 7.275 8.657 ;
      VIA 7.23 8.64 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 8.64 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 8.1 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 8.083 7.275 8.117 ;
      VIA 7.23 8.1 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 8.1 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 7.56 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.543 7.275 7.577 ;
      VIA 7.23 7.56 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 7.56 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 7.02 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 7.003 7.275 7.037 ;
      VIA 7.23 7.02 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 7.02 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 6.48 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 6.463 7.275 6.497 ;
      VIA 7.23 6.48 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 6.48 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 5.94 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.923 7.275 5.957 ;
      VIA 7.23 5.94 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 5.94 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 5.4 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 5.383 7.275 5.417 ;
      VIA 7.23 5.4 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 5.4 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 4.86 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.843 7.275 4.877 ;
      VIA 7.23 4.86 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 4.86 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 4.32 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 4.303 7.275 4.337 ;
      VIA 7.23 4.32 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 4.32 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 3.78 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.763 7.275 3.797 ;
      VIA 7.23 3.78 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 3.78 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 3.24 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 3.223 7.275 3.257 ;
      VIA 7.23 3.24 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 3.24 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 2.7 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.683 7.275 2.717 ;
      VIA 7.23 2.7 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 2.7 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 2.16 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 2.143 7.275 2.177 ;
      VIA 7.23 2.16 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 2.16 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 1.62 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.603 7.275 1.637 ;
      VIA 7.23 1.62 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 1.62 pe_5_2_VIA23_1_3_36_36 ;
      VIA 7.23 1.08 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  7.185 1.063 7.275 1.097 ;
      VIA 7.23 1.08 pe_5_2_VIA34_1_2_58_52 ;
      VIA 7.23 1.08 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 11.34 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 11.323 1.371 11.357 ;
      VIA 1.326 11.34 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 11.34 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 10.8 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.783 1.371 10.817 ;
      VIA 1.326 10.8 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 10.8 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 10.26 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 10.243 1.371 10.277 ;
      VIA 1.326 10.26 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 10.26 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 9.72 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.703 1.371 9.737 ;
      VIA 1.326 9.72 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 9.72 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 9.18 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 9.163 1.371 9.197 ;
      VIA 1.326 9.18 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 9.18 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 8.64 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.623 1.371 8.657 ;
      VIA 1.326 8.64 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 8.64 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 8.1 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 8.083 1.371 8.117 ;
      VIA 1.326 8.1 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 8.1 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 7.56 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.543 1.371 7.577 ;
      VIA 1.326 7.56 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 7.56 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 7.02 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 7.003 1.371 7.037 ;
      VIA 1.326 7.02 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 7.02 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 6.48 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 6.463 1.371 6.497 ;
      VIA 1.326 6.48 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 6.48 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 5.94 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.923 1.371 5.957 ;
      VIA 1.326 5.94 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 5.94 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 5.4 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 5.383 1.371 5.417 ;
      VIA 1.326 5.4 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 5.4 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 4.86 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.843 1.371 4.877 ;
      VIA 1.326 4.86 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 4.86 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 4.32 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 4.303 1.371 4.337 ;
      VIA 1.326 4.32 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 4.32 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 3.78 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.763 1.371 3.797 ;
      VIA 1.326 3.78 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 3.78 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 3.24 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 3.223 1.371 3.257 ;
      VIA 1.326 3.24 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 3.24 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 2.7 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.683 1.371 2.717 ;
      VIA 1.326 2.7 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 2.7 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 2.16 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 2.143 1.371 2.177 ;
      VIA 1.326 2.16 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 2.16 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 1.62 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.603 1.371 1.637 ;
      VIA 1.326 1.62 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 1.62 pe_5_2_VIA23_1_3_36_36 ;
      VIA 1.326 1.08 pe_5_2_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  1.281 1.063 1.371 1.097 ;
      VIA 1.326 1.08 pe_5_2_VIA34_1_2_58_52 ;
      VIA 1.326 1.08 pe_5_2_VIA23_1_3_36_36 ;
      VIA 6.372 11.34 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 10.8 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 10.26 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 9.72 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 9.18 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 8.64 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 8.1 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 7.56 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 7.02 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 6.48 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 5.94 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 5.4 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 4.86 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 4.32 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 3.78 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 3.24 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 2.7 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 2.16 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 1.62 pe_5_2_via1_2_10692_18_1_297_36_36 ;
      VIA 6.372 1.08 pe_5_2_via1_2_10692_18_1_297_36_36 ;
    END
  END VSS
  PIN array_array_6632d_d[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.704 12.653 4.728 12.737 ;
    END
  END array_array_6632d_d[0]
  PIN array_array_6632d_d[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.816 12.737 6.84 ;
    END
  END array_array_6632d_d[10]
  PIN array_array_6632d_d[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.664 12.737 5.688 ;
    END
  END array_array_6632d_d[11]
  PIN array_array_6632d_d[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.608 12.737 4.632 ;
    END
  END array_array_6632d_d[12]
  PIN array_array_6632d_d[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.416 12.737 4.44 ;
    END
  END array_array_6632d_d[13]
  PIN array_array_6632d_d[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.744 12.737 3.768 ;
    END
  END array_array_6632d_d[14]
  PIN array_array_6632d_d[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.12 0 9.144 0.084 ;
    END
  END array_array_6632d_d[15]
  PIN array_array_6632d_d[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.6 0 9.624 0.084 ;
    END
  END array_array_6632d_d[16]
  PIN array_array_6632d_d[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.072 12.737 3.096 ;
    END
  END array_array_6632d_d[17]
  PIN array_array_6632d_d[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 2.784 12.737 2.808 ;
    END
  END array_array_6632d_d[18]
  PIN array_array_6632d_d[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 2.976 12.737 3 ;
    END
  END array_array_6632d_d[19]
  PIN array_array_6632d_d[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.896 12.653 4.92 12.737 ;
    END
  END array_array_6632d_d[1]
  PIN array_array_6632d_d[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.032 12.737 4.056 ;
    END
  END array_array_6632d_d[20]
  PIN array_array_6632d_d[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.32 12.737 4.344 ;
    END
  END array_array_6632d_d[21]
  PIN array_array_6632d_d[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.224 12.737 4.248 ;
    END
  END array_array_6632d_d[22]
  PIN array_array_6632d_d[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.8 12.737 4.824 ;
    END
  END array_array_6632d_d[23]
  PIN array_array_6632d_d[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.184 12.737 5.208 ;
    END
  END array_array_6632d_d[24]
  PIN array_array_6632d_d[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.088 12.737 5.112 ;
    END
  END array_array_6632d_d[25]
  PIN array_array_6632d_d[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.432 12.737 6.456 ;
    END
  END array_array_6632d_d[26]
  PIN array_array_6632d_d[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.144 12.737 6.168 ;
    END
  END array_array_6632d_d[27]
  PIN array_array_6632d_d[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.048 12.737 6.072 ;
    END
  END array_array_6632d_d[28]
  PIN array_array_6632d_d[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.376 12.737 5.4 ;
    END
  END array_array_6632d_d[29]
  PIN array_array_6632d_d[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.048 12.653 6.072 12.737 ;
    END
  END array_array_6632d_d[2]
  PIN array_array_6632d_d[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.336 12.737 6.36 ;
    END
  END array_array_6632d_d[30]
  PIN array_array_6632d_d[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.528 12.737 6.552 ;
    END
  END array_array_6632d_d[31]
  PIN array_array_6632d_d[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.008 12.653 7.032 12.737 ;
    END
  END array_array_6632d_d[3]
  PIN array_array_6632d_d[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.584 12.653 7.608 12.737 ;
    END
  END array_array_6632d_d[4]
  PIN array_array_6632d_d[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.16 12.653 8.184 12.737 ;
    END
  END array_array_6632d_d[5]
  PIN array_array_6632d_d[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.448 12.653 8.472 12.737 ;
    END
  END array_array_6632d_d[6]
  PIN array_array_6632d_d[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 8.544 12.737 8.568 ;
    END
  END array_array_6632d_d[7]
  PIN array_array_6632d_d[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 7.872 12.737 7.896 ;
    END
  END array_array_6632d_d[8]
  PIN array_array_6632d_d[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 7.104 12.737 7.128 ;
    END
  END array_array_6632d_d[9]
  PIN array_array_6632d_q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.512 12.653 4.536 12.737 ;
    END
  END array_array_6632d_q[0]
  PIN array_array_6632d_q[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.72 12.737 6.744 ;
    END
  END array_array_6632d_q[10]
  PIN array_array_6632d_q[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.472 12.737 5.496 ;
    END
  END array_array_6632d_q[11]
  PIN array_array_6632d_q[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.704 12.737 4.728 ;
    END
  END array_array_6632d_q[12]
  PIN array_array_6632d_q[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.544 0 8.568 0.084 ;
    END
  END array_array_6632d_q[13]
  PIN array_array_6632d_q[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.448 0 8.472 0.084 ;
    END
  END array_array_6632d_q[14]
  PIN array_array_6632d_q[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.64 0 8.664 0.084 ;
    END
  END array_array_6632d_q[15]
  PIN array_array_6632d_q[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.408 0 9.432 0.084 ;
    END
  END array_array_6632d_q[16]
  PIN array_array_6632d_q[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.264 12.737 3.288 ;
    END
  END array_array_6632d_q[17]
  PIN array_array_6632d_q[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.168 12.737 3.192 ;
    END
  END array_array_6632d_q[18]
  PIN array_array_6632d_q[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 2.88 12.737 2.904 ;
    END
  END array_array_6632d_q[19]
  PIN array_array_6632d_q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.8 12.653 4.824 12.737 ;
    END
  END array_array_6632d_q[1]
  PIN array_array_6632d_q[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.84 12.737 3.864 ;
    END
  END array_array_6632d_q[20]
  PIN array_array_6632d_q[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 3.936 12.737 3.96 ;
    END
  END array_array_6632d_q[21]
  PIN array_array_6632d_q[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.128 12.737 4.152 ;
    END
  END array_array_6632d_q[22]
  PIN array_array_6632d_q[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.992 12.737 5.016 ;
    END
  END array_array_6632d_q[23]
  PIN array_array_6632d_q[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.28 12.737 5.304 ;
    END
  END array_array_6632d_q[24]
  PIN array_array_6632d_q[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 4.896 12.737 4.92 ;
    END
  END array_array_6632d_q[25]
  PIN array_array_6632d_q[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.568 12.737 5.592 ;
    END
  END array_array_6632d_q[26]
  PIN array_array_6632d_q[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.952 12.737 5.976 ;
    END
  END array_array_6632d_q[27]
  PIN array_array_6632d_q[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.856 12.737 5.88 ;
    END
  END array_array_6632d_q[28]
  PIN array_array_6632d_q[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 5.76 12.737 5.784 ;
    END
  END array_array_6632d_q[29]
  PIN array_array_6632d_q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  5.856 12.653 5.88 12.737 ;
    END
  END array_array_6632d_q[2]
  PIN array_array_6632d_q[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.24 12.737 6.264 ;
    END
  END array_array_6632d_q[30]
  PIN array_array_6632d_q[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.624 12.737 6.648 ;
    END
  END array_array_6632d_q[31]
  PIN array_array_6632d_q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  6.72 12.653 6.744 12.737 ;
    END
  END array_array_6632d_q[3]
  PIN array_array_6632d_q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.296 12.653 7.32 12.737 ;
    END
  END array_array_6632d_q[4]
  PIN array_array_6632d_q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.68 12.653 7.704 12.737 ;
    END
  END array_array_6632d_q[5]
  PIN array_array_6632d_q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.968 12.653 7.992 12.737 ;
    END
  END array_array_6632d_q[6]
  PIN array_array_6632d_q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.256 12.653 8.28 12.737 ;
    END
  END array_array_6632d_q[7]
  PIN array_array_6632d_q[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 7.584 12.737 7.608 ;
    END
  END array_array_6632d_q[8]
  PIN array_array_6632d_q[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 6.912 12.737 6.936 ;
    END
  END array_array_6632d_q[9]
  PIN array_array_6632d_w
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 9.408 12.737 9.432 ;
    END
  END array_array_6632d_w
  PIN array_array_6632d_widx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.504 12.653 9.528 12.737 ;
    END
  END array_array_6632d_widx
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.672 0 0.696 0.084 ;
    END
  END clk
  PIN counter_delta_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.768 0 0.792 0.084 ;
    END
  END counter_delta_ready
  PIN counter_pop_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 8.736 12.737 8.76 ;
    END
  END counter_pop_ready
  PIN counter_pop_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 9.024 12.737 9.048 ;
    END
  END counter_pop_valid
  PIN expose_executed
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 9.216 12.737 9.24 ;
    END
  END expose_executed
  PIN fifo_north_pop_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.416 12.653 4.44 12.737 ;
    END
  END fifo_north_pop_data[0]
  PIN fifo_north_pop_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.272 0.084 10.296 ;
    END
  END fifo_north_pop_data[1]
  PIN fifo_north_pop_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.6 0.084 9.624 ;
    END
  END fifo_north_pop_data[2]
  PIN fifo_north_pop_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.216 0.084 9.24 ;
    END
  END fifo_north_pop_data[3]
  PIN fifo_north_pop_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.448 0.084 8.472 ;
    END
  END fifo_north_pop_data[4]
  PIN fifo_north_pop_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.488 0.084 7.512 ;
    END
  END fifo_north_pop_data[5]
  PIN fifo_north_pop_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 6.912 0.084 6.936 ;
    END
  END fifo_north_pop_data[6]
  PIN fifo_north_pop_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.88 0.084 2.904 ;
    END
  END fifo_north_pop_data[7]
  PIN fifo_north_pop_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 8.928 12.737 8.952 ;
    END
  END fifo_north_pop_ready
  PIN fifo_north_pop_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.864 0 0.888 0.084 ;
    END
  END fifo_north_pop_valid
  PIN fifo_pe_5_3_west_push_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.648 12.653 3.672 12.737 ;
    END
  END fifo_pe_5_3_west_push_data[0]
  PIN fifo_pe_5_3_west_push_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.168 12.653 3.192 12.737 ;
    END
  END fifo_pe_5_3_west_push_data[1]
  PIN fifo_pe_5_3_west_push_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.696 0.084 9.72 ;
    END
  END fifo_pe_5_3_west_push_data[2]
  PIN fifo_pe_5_3_west_push_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 5.376 0.084 5.4 ;
    END
  END fifo_pe_5_3_west_push_data[3]
  PIN fifo_pe_5_3_west_push_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 4.032 0.084 4.056 ;
    END
  END fifo_pe_5_3_west_push_data[4]
  PIN fifo_pe_5_3_west_push_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 3.552 0.084 3.576 ;
    END
  END fifo_pe_5_3_west_push_data[5]
  PIN fifo_pe_5_3_west_push_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  2.976 0 3 0.084 ;
    END
  END fifo_pe_5_3_west_push_data[6]
  PIN fifo_pe_5_3_west_push_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.36 0 3.384 0.084 ;
    END
  END fifo_pe_5_3_west_push_data[7]
  PIN fifo_pe_5_3_west_push_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  0.96 0 0.984 0.084 ;
    END
  END fifo_pe_5_3_west_push_ready
  PIN fifo_pe_5_3_west_push_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 9.12 12.737 9.144 ;
    END
  END fifo_pe_5_3_west_push_valid
  PIN fifo_pe_6_2_north_push_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  4.608 12.653 4.632 12.737 ;
    END
  END fifo_pe_6_2_north_push_data[0]
  PIN fifo_pe_6_2_north_push_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 5.472 0.084 5.496 ;
    END
  END fifo_pe_6_2_north_push_data[1]
  PIN fifo_pe_6_2_north_push_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 5.088 0.084 5.112 ;
    END
  END fifo_pe_6_2_north_push_data[2]
  PIN fifo_pe_6_2_north_push_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 4.704 0.084 4.728 ;
    END
  END fifo_pe_6_2_north_push_data[3]
  PIN fifo_pe_6_2_north_push_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.648 0 3.672 0.084 ;
    END
  END fifo_pe_6_2_north_push_data[4]
  PIN fifo_pe_6_2_north_push_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.456 0 3.48 0.084 ;
    END
  END fifo_pe_6_2_north_push_data[5]
  PIN fifo_pe_6_2_north_push_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  3.552 0 3.576 0.084 ;
    END
  END fifo_pe_6_2_north_push_data[6]
  PIN fifo_pe_6_2_north_push_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 2.784 0.084 2.808 ;
    END
  END fifo_pe_6_2_north_push_data[7]
  PIN fifo_pe_6_2_north_push_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.056 0 1.08 0.084 ;
    END
  END fifo_pe_6_2_north_push_ready
  PIN fifo_pe_6_2_north_push_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 8.64 12.737 8.664 ;
    END
  END fifo_pe_6_2_north_push_valid
  PIN fifo_west_pop_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.56 0.084 10.584 ;
    END
  END fifo_west_pop_data[0]
  PIN fifo_west_pop_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.176 0.084 10.2 ;
    END
  END fifo_west_pop_data[1]
  PIN fifo_west_pop_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.888 0.084 9.912 ;
    END
  END fifo_west_pop_data[2]
  PIN fifo_west_pop_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 9.12 0.084 9.144 ;
    END
  END fifo_west_pop_data[3]
  PIN fifo_west_pop_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.832 0.084 8.856 ;
    END
  END fifo_west_pop_data[4]
  PIN fifo_west_pop_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 8.064 0.084 8.088 ;
    END
  END fifo_west_pop_data[5]
  PIN fifo_west_pop_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 7.392 0.084 7.416 ;
    END
  END fifo_west_pop_data[6]
  PIN fifo_west_pop_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 6.432 0.084 6.456 ;
    END
  END fifo_west_pop_data[7]
  PIN fifo_west_pop_ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 9.312 12.737 9.336 ;
    END
  END fifo_west_pop_ready
  PIN fifo_west_pop_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.152 0 1.176 0.084 ;
    END
  END fifo_west_pop_valid
  PIN pe_5_3_counter_delta[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  12.653 8.832 12.737 8.856 ;
    END
  END pe_5_3_counter_delta[0]
  PIN pe_5_3_counter_delta[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.176 12.653 10.2 12.737 ;
    END
  END pe_5_3_counter_delta[1]
  PIN pe_5_3_counter_delta[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.792 12.653 9.816 12.737 ;
    END
  END pe_5_3_counter_delta[2]
  PIN pe_5_3_counter_delta[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.888 12.653 9.912 12.737 ;
    END
  END pe_5_3_counter_delta[3]
  PIN pe_5_3_counter_delta[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.6 12.653 9.624 12.737 ;
    END
  END pe_5_3_counter_delta[4]
  PIN pe_5_3_counter_delta[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.696 12.653 9.72 12.737 ;
    END
  END pe_5_3_counter_delta[5]
  PIN pe_5_3_counter_delta[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.984 12.653 10.008 12.737 ;
    END
  END pe_5_3_counter_delta[6]
  PIN pe_5_3_counter_delta[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.08 12.653 10.104 12.737 ;
    END
  END pe_5_3_counter_delta[7]
  PIN pe_5_3_counter_delta_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.248 0 1.272 0.084 ;
    END
  END pe_5_3_counter_delta_ready
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  1.344 0 1.368 0.084 ;
    END
  END rst_n
  OBS
    LAYER M1 ;
     RECT  0 0 12.737 12.737 ;
    LAYER M2 ;
     RECT  0 0 12.737 12.737 ;
    LAYER M3 ;
     RECT  0 0 12.737 12.737 ;
    LAYER M4 ;
     RECT  0 0 12.737 12.737 ;
    LAYER M5 ;
     RECT  0 0 12.737 12.737 ;
    LAYER M6 ;
     RECT  0 0 12.737 12.737 ;
  END
END pe_5_2
END LIBRARY
